BZh91AY&SY�%VJ 1߀Rx����������`7}۽�k��'N�A�T4M��I6����L�� ��4A$I�&�&�dz��  �  �)�cD4   � �� h�   �2d�b`ɂd ф``$Bz&4J~MSjzji�jy �SF���������X��q�BD�Ւ�� �n��K�G�j�1$�E��r��`
��.�i��lE����¦�4	���J����+f����ZG#I4�%�8��FuIa�z��@LZ��l�"gj�$f���G(fR��g�m+��҃]�H�S�MԾ�O��1�\7R�N�`e�[\4� ܼ��I�t�U�ٵ,��y�`x���.��|����4u�(�7��M&9bg!���;�Q_q�� ���3�D2�
�t"��lQEa���r+�b
��Q5-�4�D�a���(�Rt�3-�Y�Y��me,\�'#�ɜD�"l�����l�@���gړ!Hh`���ɟ!�<�,��r��)�h��'�N�EnUv�AjC) 
�)@D:�\VA$�I�&+��1�
�*2����w��&l�����wY;���ߗJƗ�����R8O��^5V��ę������[0Y�.T�.���&���ϖ���%�1�hq>L��-����hc6$�����S\��_��ඐag�����]�(%���	;E�yׄw��l�c�X�؞j��M%����a��3l�����/tsH��Dwom�L�Z +��p�2�
j�)_']A��i���U�z:TD9{��G.H���ַV�4tkΧAR�JIp��M��KU`:f�i� ���i�ƛP9�cR�O�9H,n��a�:�:rU����L�aYC"e���$��~^�k����D��((�H�p��+=:�ύF����JE�PWy�cd�	k�]5f��F��c"�S�O��(8LS��(�վZ�Ê���±� P�}�A�!2�S$Cpm?tA�L��4�1�����7�\T���+L�-%q�:�f�mh�ji��w�i^�6u��Er*C�.��V�(1]u����Li��8���T$0i]6I$LEA�N� `�8c!��[PAր�,��U���HbR�-����-j��!�
��մ���鋁����wG2�ٱ%���0Ϗ���� <I{P1�b�F7ߤ�j�Y�9��[��_Z\���Af¹/���`(;_��_"���a��O�2�I�8J�ؓ8�D�j�<2??y��5T\s���`
���&�G%����d�2�k��	�EM����(0l��n�T`�RR1��2�hǘ�ݟ#$�uٙ�<�vd$Q.������-�W9ƅf�.kg�B��U��$���_���sA�My�!#Z�M�	��v[#iYT�*#R	�.'88ȆdT�-��c�u��A�!�y�<JЧg�����H�
��@