BZh91AY&SY��: _�Px����߰����P8�7LEBQ$��LFڦj0M4i�h�d�G���5�F��I���d�  �'��ji24��2h�����9�14L�2da0M4����$�OSh�bF���224   �(�"T��_
 ���eI6��P�cIv�V�Z�����sd>S9ǋ��2���u'�sl�2H\WL]yFST����j h�<bINV���\�^cs3�1�����B���)�poyA|�T}�EmZ����k�({M�7\���o�	�/�uOEl����׮M5m����d�ӹ��3�ū��]�(q��椔n��r��VD��3�у$��&��*R�VV��13g��k����)8����|'�t�H	����e�{K
��E��٥@�p�N�^�=�>�$�Î��i�����PL��A���Da"u\YR�׉G)}�ί�R(�	�!�Wpp����Q��(O�j��O�ꧦ�G���r��R�&��C�O�ݶ8c
8���4Ӧ����.U,k~��	�4��QL��O�N�,B�����>\	����2A�v���N��v*"lP��-]�΅�^b�vūi��'v-P���XK��6m�k^�
�*�&�+Xօ/��'�@�\p�F�8}i'~�J��t��YU.�h��$�"���e��J���<kTXG �P����>�%"��@��T�`�X#}�ؠ��t�z��+� @L+N��������8w�l���Ģ�ŷ[��_�o���dI-^5WC�Dh�琥����B��Vъ�����1�u����ߠ��)�Ȥ�