BZh91AY&SY�P{- _�Px����߰����P8��b��BR*yF���=CCOP�M0@��COP1A2&�i��!� ��F��� h	�j��dh��F� F�Ph4d���`F�b0L�`��SM��	4�L���   4_I�!��Z�R�пl���M�g�P�kIs�cJƭk�����H����K�e֐5�צ�v�ٞ���N�)L�3m�-�P��*�%'r�Xf{����2����c���`)�(���K�j�*����%���%�z�S�z��_�
�&��߇6zn����''�hci��l��}㠹_oA
n��)��VW}�[Q�[��F��.=��vёA�sC3�Mb�^"�<g�T�v��{~���H�O�,�-�C��ޮ5l~���!CU8�񉒍����Վe��e�iru%Z�ņ�-�I�eI�dK���EF��F��F��A�!�T}�)�)�1ȁI,+����}�n@������Ź'cD�=z�NՌ(�H񡦝f�\L��ah]f[���'0ҧ��׼�17�(����[�;u�E�����\�����q�T=ڡX�~}�t�2���V1ңB.@�#�T0c߼�^4�Y������T����)^6#L�� ��I՘�R���76@֋�m$R��S��Y�=��7	 v�a��zi�*��gޅ�� h���oga��8��c/�&��9����^��� @Ʌi����%[������4Dp������&�a����dIm^����Da�"2O)S"�	������E�!J��@چ�Yȇ���)����h