BZh91AY&SYbym _�Px����߰����P8�7N��j��H2` M	�4� 4 m@�&��B ��M   ���D�����)��SOP hP=@�101��&$�5M�jz4&�4��4   �=BD �+��A�/�&��I���	i-�Q�F��k:�:�D}%-Q��z�eH��r塶e�D�ҹ"�e�Ԗ�M�;�T�%Q�9��������)�F,���;���������3Os{�j��
8���;��<�PI����t�J�c�Y�e-�'~����b�ӫm�j�w�����P�TGnr&�>��0b�M��E��	R ��܆5j�RNvkl;��x�x<M�-�(z�
��m��$���T��y�1�*^��9��R��8@|��)����Y���IZ>K-	��-`~���eDa�#�]i.g�d�|��|_��V�?j��q`A`>��t�/9���(ߡ�b��᚞�j5jx 6��i�|aF��rֆ�s�*�Rٲ�B�]z<�$�&�=ex���"��+�;��,p�֑����<���Ŵ6O��=�1�%U�˿��.
���jPRa�]yQ�u�[!X`4)FRk�	1f�p:5�W;����d��Ąa"1d.�t�d#�%4�l�l���KuQiEe�,L���2"��Ï! ���Bԫ��n~�3� �i�d�)+�Z�K^.!%(c�9�f��t�W�ɏFdɁ0��Q �i�e���Z�_LmyT���5͕/�Jʝ�K�&B��	M�����J��+�M���&ъ�Yg�cb��`]��ܑN$؞[@