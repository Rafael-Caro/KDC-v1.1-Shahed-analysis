BZh91AY&SY��_� <_�Rx����������`?zۜ�3�Z 
�"j����=F� �@�@A$��ɐQ$�M 4�������0L@0	�h�h`ba��B��=#M��hш�  � �`�2��H�h�������y4��2M4d����Pr���b�4��%���I7������9��#" BV#���IВ��#��6��6�S����|�X�V���b �ʬ���x*�K�J�J$��	����{Y劸T�j�{�=^�h���~Ee:�3��x�gf4p�x�Q�o ��C�Jq�ܟ����+K΁��!�����$
�7����K�����$�e�0�L<�_}0�c9j��~7u�*�7��$>m��$ϐag��g��ol�X��D��_���K1���%��+�)�D��	 �����U��ǔ�c�Vғjk5���Vc8����Tm�4ĥ��d��6k���޾ĿK�k@��� ` .8�8�5����'Dr�a�Ŝ��V��K�����T�'x2i�M%5uz��rB�ə�EĲ��xe)1�7
(2��@`����fO� f+G,\�Z���8u��T�R�5�W�6��;D��-��t�&!gP�ui�f�H85�\=uc ִ1����Ԟ����@ءU�eˇ��oE��s+�x�?�����������Eڂ�]�B$wi������*;mz��S(SG�c/��L���6�� ��x��9$L{�:��٦EW@[�vD��)�ؤ}��M������G�y�Ġ�ɩ�����`���_Ke��i����曽��b\J��X�,B�]�A �iV�q`��[۔���J�}��$q�Y$����~Z�4l-*bL����j��a��f��b=+�
�:�e�bg�a�v�������;� �A��2T�V��h�i)�O��	&)�xH��vG�b�5�3��A�@�-c����y�k��y?Er�p��t5�ݸ���?<�1���(�w���L�����	s�xh4�P:����E�,è0����*1�]vCAUj�&4�1!�$Fb�ge�C�%Ɔ�I`At'H `�8c!���h������P�	Hd�4��r��Jl��
���\Tݿ�V�0B{�.�~��EѳbKUm�0˟�w����"G��ٱd#Fl�MF�a5�Ð�������K�3��96�{�x��{�����:|���<�"x'	A����rC����D�H��ݖ,�
"�JƚsI�'�gAbNJ��\���s��]�hpsޜTX"o�D�u��POO,3��1����p���2֌����)K���;zGD�TWGD�S(i��� �)P�ǜ��[[��&���8��jEv�&#!Х�6�� �b�F���n��dR�����o�g��R{�:biG�ȵ
t�Fo�]��BBf�~�