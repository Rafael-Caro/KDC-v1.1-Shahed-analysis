BZh91AY&SY�{�  �_�Px����߰����P8�7N�j��H2ƞ�� 4��DѠ @�&�M��i���F�hi��M$D���`I��M  ��101��&$�5���&�3B24@ �х�$BT2k�D��������P�kIt5cJƭk�ƾ!��C�>�;#{��2��5�צ��Kl�Y$.-��Q�)\�΄D�|�I)��f�<mh7��*Q��^x�,U��T"_�S��]E(�6�QTHP����]!5<X\�_s��|4�Ō��Vp���'&�����km�m�;�W��t�������$�uW�e~�CV���a�a�(o�Ll�.j�C�G)7C4�=�Z�2�ɵ�&�D{��^�c��E2���D,�hmM`����9�Uc��ZL�A+�SD�h��PI��!'�i��70?Phd�(�3����'��z�,�~�K�"�CP��x� �!T
�rmVR�����#�g�T���$�h�Ƽ�F� s�4�Z�g���Э���')8�*8�Sn����b�.�o2�-٬�
0y�C$�e���	:�\RP�	Ȅ�%�u­-�cR����j��m"��Z�`.�PK��	X��q�kq���`�5Qp��F2FCL���D�I���R�v�5l��%�j.,U���!�X�=����� k����4J�T�q����8�5���x�[���\"
P�fr	�f|AA;�:���D���G���^f���R}Z�l:��R(�6t�I;/:S��f1�[�-S��p�&�R�S[w��ђ���[�1�s3p�E��H�
 �/w@