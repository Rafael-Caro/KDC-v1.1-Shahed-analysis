BZh91AY&SY�5  �_�Px����߰����P8�i�vn��(P�D�==D���!���4h@@������jh0��!�i�A�z�H�HL��&�hi6�  �=C@���&L�20�&�db``I�5OS`Pa�4     _)�!AZ���B��ZI6Oȡ"ƒ�j�*�c\��1��z��ҕ��C��l k��)M�M�(P.,���Y�i/��m��hJ�E""Z/Xc��e�rq��QvCN���X,���E�����/�8��&r�>���&��)66MTi�i	���S�|�ަ��N噍�km�l�E���]D(q��#�4%�,�������!�����(aXʖ�(X�r�y�Dv?H�|�$k5�U�Z�.��f�+�ݡ�����t���7��f�-��+ZB�|+�$�u��<y|�1:y,ә*���F����.5ғe��=O��~�K���C�W��X�X�%�Δ'�u�J���ςX�u��E��9��
L���Q�Q�P:lCM9�,qJrrT�-�K���>i$ �d��ڛ(�-�T����c�D}�P�<�e�N��$�$�\���PD��^��*HW-)��<?�#�A&�ņ'�qJ`	��[��=����j�6�mE�1!P�F���FP��cD�;.���5��s؈���zdA֤G|�D�ǮJ]`e�::Kv�6�r:@�q�ф�4�ۚ{�Z7��`��+�a_�����cЉ D�R8@|W��:{�&���-$ �7���P��B�SQ4���KG	A���C�^@r�0NWW)E�B�֭�62޷�cb�̀dʋ��H�
1�f�