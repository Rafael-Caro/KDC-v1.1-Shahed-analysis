BZh91AY&SYA簓 ;_�Rx����������`?z���!�U �2�L����L�F��2�� i��hi�     4  �=S�i���hL�2a4  zH(���Q����چ0& � q�&LF& L�&@F �"@�	�`Jy�➛ByL� 4�52m&T?�	Aւ���i.!KsK�HI7����W���d@��G�%�'�J��D���Ŷ"���b��(�v�
�
��ij��&�"�lY����� �����#6ߘ�q�tz/��֊`��:�0�K��mK��4��w�1���V� '(�,,��3M�U�9yV���i]>8]P��8̕R@��	�4I%�z0����.�����������0c���|����.�7ï� եA���	=�~%�MN�Sߕ��Q�5�"C����ث�s3kEIۅ*�S�!;�M����J�T�l(�y����WV��a�b1�T�)��[�C3��RY����/��^tY[B ݈�C[{�^�q8F��$0W��#@�l�Q{�߲�U%���qi8pKH�LBJU�&�ɤ�\'X%�oZ�V�<-1U��XiTa�a%��bbh `�NN������>��)6���M_��{
j���x�=f:�h��R�Y+𦛥d�!/-��>3�sL��$��e�b���������0x��^kb�X��7����A����g���/z�{�b$|���i��.;� �O��(SG굗��sMa�f� }��QyGT���G�F�6ȱ�
�0�h��5����ƙ$D��+//k���9�()I����C2F;忻r�gBsQƝkv�K<��^\J�pOm�[L�]� �D4�+��W"h�[R��ˆ̶���H��P�(�2+Ӗ�͜
�5&[b�Iux}��T�m_�3$�1AU4��_�&��o?:�W��T��A\�k$H9/`���[����EIO�~w$\$vLS��.���}a�I��s��B�iBi�	��.b2�m�<���^cLlhc���Ø?�"��ol�5��,������U3�Ga�����m_ 8z���"�(��2��L\��jz��Ƃ�t��L�&D�f@3-A!�H��D�P ��0s1���B�� �Y�TD���&BR)M-��Gю%65
����)"!�˧�+1>�YH�m�[�]&�~���}��y>�cg�F���N'b�è�5 �NRnD$�
R��t�
�������v6�I��I"y'	A�	3�$U����C�n����a�h
�,��i�&L���b�9*�,��#6[�M��������WF2l�J)CEU%#`�i���;�DDff��ɷ�/���*���F�6�g����s9��Qbdn�uT�&��H�,����bh?t׬��7��\��C�ldq*`�q��7(���c�k6��5׎?7I� �� ڏ\�T)�ۈ�����)�=��