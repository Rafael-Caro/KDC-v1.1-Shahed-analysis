BZh91AY&SY;�{  �߀Px����߰����P9�0�%��JB�OH�y#@����L�COP%�b$Ɍ�h�� �� " ��?SP�=�<�@  P�0&&�	�&L�&	����jMM�A��@    TO�H�hb��"0��eI6Oȡ"ƒ�5V�Z��\��1ɐ����8=/b��aSk�[T�uÂD.4�=E$Q��c�6��3	DY��1�:�>�&J"�Wg���B�^��a$hriyٗI4ow)[@���fT��rR�`�j>r�=G=M
���AA�������6h�\lm;�m�3-�t�_�y
p�ڤ�wşw5��n�b��É�p�L+ 5I6�J��u����5���KFe�����>���.�\�tx��6�3���-�"�v;�u0�3��ȅ��L�a"��=K�b�2g�Ph|��eH��jOcG(ؿ�W�(�J ��u
v�
}>y�Δ'�\�<��ߣ�Z��\���S͚$��O;�����@�Zi����͕,k7s�I !Y&,6����*�4�_X	�>��E�a��YI֠d����
A�eK*U��R��⥚xN����H~қ�a�iM�3����Zx6��3-f���o9�֢���$�F�(}f'�J��t��Y��q*�x&De��z41���,l#��T��e�5��$'<� 0�Z�ܞ�0�����"�p�+���?s}�bD�(�E\,.P�~ܳ��F�iJ�ƛ�t��34꬘��KG	A���C�\@r�/�WW)E� ���h�R�[�y�6.vk�ȷ�.�p� w��