BZh91AY&SY��� 2߀Rx����������`?z��=�L�� ��^�E<S�H2h'�M=�&� l�h�� i�  @  iO�I<�L����4�  4 )�	I�OTzi=M���h�1���9�#� �&���0F&"M!�14���z��"yM4 �ɓ+���Ac�b�D��KcK�H��~o�zB?j6�BIQ֢P}�u�q@FC �g��~^����asE�#��d5h�q��8re����lF��mԦh�619�C�d���k]ࢴ�8�E���=3	�Y�/l)|�A�		��C���v��*�W�c<�D��E�3�Xa$�WT�I4mI�5$߽3�:�.v8 ���V�t� !�R����Ph��3���T�a>�����W��H�u8�8,U�8b�A�o\(,
�Bv�QR�3$�G��䱬C� e�����V�6r A�8M2��V,�PCŧw|?G�$#&�$�I$y��D�.��q�ǚE���L���=��G%%�x*K�0�����'X�ɀNu���W���*�U�ƕF��jjz�!W��)�#�:���3?.�	����)��������4�>�B�n�
��uA���Pm}�6��� \��.�c �\���9�&
8o@76yO	�\�D]�aU��E���g�Hp��XKq��	zE��y��z>f��ڈ<ޯ�
������scN!��� y��b�G4�DG�5�y�
�0�h��E��_��)+t޽�v�ҫ��D&VR����aESU�i��Q�U;\��]��k=ؼ��4�J���^���B��	C
ٝ������i��e�+�_o(97I9f�$v�῝3Vҥ���]�J\��"�*C5��4�ؠ��F�/�&w�9��u��U��u&WPWA�1�B	��.WoW�{�5IRi�N�(�IƂ���d��v�8����]�� ��8�#�-�.�3ŏ��/�m��1�`�y���_@?�"�S��q3�Ĝ����!�j�������e�ֽ 4m�0.!���;)4�`�ņ#3��p�4U[%�4��H�F��ie�C�+��R("��+��І�3���]W"p��(BR2f�k��8�3�,��� ��;t���T!F� �F�����nFK@���=^�j3�I�56��5hѬ�l�&��y��L[��^4��KIu_������i��4s���җ���9|�"�'	A�RgT$HQV�3��qFˌ���KH*�^�J�i����!���.�"���d[J��#_�ƑYȺ��PuƕU*MC�z�m~<�p�-��	��xv��"���]*���aB�f,L���j��#I;l/��}M�5�$�s�-��A�y~2n*`�a��6�-۠7�o/��U���p��d�q-� j ��W!�.�p� ��