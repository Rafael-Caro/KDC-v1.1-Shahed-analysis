BZh91AY&SY�f�D  �߀Px����߰����P8�=�V�Q �51���4�m	�� ���OCHɈQ�h�hL� 	�i�F�2)�b�d@z�������a2dɑ��4�# C ���ѣ       Ɖ�!A^��QF�_�(��I����BE�%��ZUj�d�@�I{��wG����}�?h����9)$���-�F`5RWL�Z/X+�����tM�c���vV���N?����&�{�s5F��3_q���9��
4Z"���m҈���1����" ��aդ������}�SNͶ���;Qz�~]�\��x��uRJ^E��/�?�0�6�Oh��Zx�U�9Iu3Cc�5��,���� 3Ů>����g����%��0D�.�)&(Y�%�@�잠:
n��U�wf��/�f*M�yq֙��k��O�DabZ�])6X#��g��~
OR!�5
�W�2@�'�Y�Ow���1k_o5��5)�I!�O{��65�m�M�i�Ms��~z���vq'@ң�E7m�O��W�Y�������O���C$|JcIH'����tdY�H�
R#ՠKIu6��K�	��!6[E��Z��
��PI�7��3v�Z��Up:�E�fB4I�2��d2O��9J��i���*�MȱU}�pM+���c�aP��:�����f�o�̯+�#�Kf0)2@Ū��_r��P�+0��Lcb���d�|����X�	1$ ��F7C�R}]v���)k�2]$���т]�3�` 6���(��O����<��#�����3T���>A������$_���"�(Hf3H� 