BZh91AY&SY�X�* _�Px����߰����P8�7L�M��Q ȓтi��@m&OHhM P5I�5<� & hh $H I�&��D�D  �=C@ѓ �`A��2`�Jej��zd!���4  �|��!X����!~�6��M���(H�Inj�*5V����1��zH��Z�����ʐ5��D��Cl�<��x��ɱ�
��JnDA�@���J���2�NR�d�<T�-����
�o��$�Z�I9�}�R�$�r}mi��ID�0R����9�s�3�o��g�&f�0[4����w6� f�鼱_�y
p��r&�>��]6WI��a{&p�F�-T�)�Z�����M��kg���'@�l�!���t�nk�Ev¡5	����I�B���P�A�dθ7hVd��Mi��0vr�|�;Gx\��A��ʈ�BGƶ������������A���{g cꁒP�e��&P��T؎ZS���n��[3D�D���i�r��2i���K^�)u���%�3 Փa�uC�Y�PF�!J�Z h�>TJ�$ k��ms�Ǵ�<�UB)D���8��q}.k��ʮ����".�G���Rl
	1�}o5s��q� �b-��Db4�Z��A�d�^2Ji��X�YQ.z�Ҋ��A�j#��D�źN/\xA�J�^&.,��P�<�@0�I^b�~Z�9q�VR��h�� +8�۟��Z�"D���>ZX-!<�k�� �/bHc\�S�����n�
&�8N�[�`Õצ��Es��y�d�m�Ֆu��6-���ȳ�.�p�!��@T