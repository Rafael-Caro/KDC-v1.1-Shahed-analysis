BZh91AY&SY��d _�Px����߰����P8�0��	DC!j~��D��2h h��`LM&L�LM2100	M'�22&�4��  h4h9�14L�2da0M4����$�SSz���Bh�OH@  ��4���������!6��M���(H�Is5F��]�+�1��r#�)k����2� k��T�ש�f���r��&̅�Kk�2#jb�T�-D�ک��rI�7�>��`�W�z7B$��8vpn5ҏ�E$��(P�o��.�J�SL���P[�T��Ҭ�
Vu��|5�ǫrō�V�d��x.���B�|��țt����QY�ɯ���ׄ�) =R�"�r�R}��?G:�Ϙi�֘�l.������G���s���	5�j![�c�S	g�5�+�vY|r��)���@�Q.B��6�ő2���&�#nΔci�����?��t�lC@��cAcMR��y�y��\��4a��`t�զ�LX`�?S�Lp�
5��i���K���BԿ";���Sq���z�Ⱥ�]��U�Tgg	/2<�#$85�Ym9�
㾦<䪡�Y���r��v�,�����ص3���EI:���;�f`�NU�L��p.�y� �d\#���i��@;�(��d�ӭҳdg�\�EĔ�ıAe��5���B@B����2J�]l61�P�<�b��P�-;TSSֱ�0�Z:� +7B�S���ZN8�81@�`�ژEo0[��S�3��ﶢ$��s�B\%���1�{E��y��������WW"�����h�N��S�1�mg�E���H�
8 l�