BZh91AY&SY��� ?_�Rx����������`?zۜ��Z
��jj�M&e4h �@@�A$�����yLA�A� �hh9�#� �&���0F&�4I����&��h 4�`�1 �&	�!��L�������Ч�Q�@Ѧ��h�#FK�?�%�>LP &���$�����Rl�ߥ��~ǘ�i\}#����JJ�`��"@�g��e�Ā��|�T�F��#� �Qɱ�M�B�h�q7"@�Aòt���nm�=�bT��U(�l��.Kq� �����Բ��3J��:�x瞫F#Y��p��o;��q[H�Z����ʂ3P5h;f�]:�R�I%�rRvRݖ���L!y;+�Fq���ݛ�"�`ޭ|��1�ZD�#�K
���bZ��e�d�50��������]��;Y�}��WC�gTU����0�=�Vd�3.�̃&Qx��K�0�9���2�`��^Y�p����.u��^D � .V������m/����,�,$s_"�)9*YU��Al˫K5�e�EEeB�;���+�eJ1�,YHd�0Y�zݛ'� f2��.v-�����Q9^����^u�>���f��baB-S��Q 9-�����Ң�ѐ���������<�c���q��_�7,Hb����n$���_5�[��j�XV��g������Z
	ȳ6$H�a��=h���z+v���(SG�c/��ʅ���6M� ���"؏^��4H�Ӛ���-`��b�5�q}�6�J���q��6%UMOD���5ȷT�sҵ��Z�ܽ���dՉ�&V���-iǄ���bĠc0q!��h�ڥo��d�KcN��Y~��$s�THu���Rf���,�v�������P��5/��JA�F���5//F�3�Q�u�u@��<�l�A �yά�����$VJ}s����;�$x�Aב��k[��L���s����GSDU�<'��|�U2�h��v����qS'ǌ�1�������C/�3cGKH%Ƌف�z�h��3�"/ P�̈M��s��f�(��ɍ4��Hc���eײ�!�H��a��D�Tf��c�2 {�ju�9�2��K4�d%!����VeV8��kPE�Pۻ���\���\�x${�zN�i-4���\~�g����$zځ���B0ϟA��\&�8t��A��)r�K�����⃱������;"|���;����􆴙�$U�߉������~�ૼc�w�lT���*�x"7t��SP��t<�o���Ax��d.3w(���Z����A�*J�	��v&)��33��	$E.Mo4�i,s)"FH�Gr��XҎ�a�S�Z�9�
�Mv�4��Q#�HԤSaBb2����VfA�uhH�ٱ��F�RfAE���:'�ۄ��B���N�5�3���H�
�ܓ�