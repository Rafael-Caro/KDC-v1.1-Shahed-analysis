BZh91AY&SYʹX� <_�Rx����������`?z۸����� �I��S��S�OF�x�=&�@�L54h6��EM�Lɦ�    � 2dɈ��	�����4��SS�i224�=L�( 242dɈ��	�����$PD�M�ȏT����3J1�����L& ��؂�͊I,!K6�֐�o9���W�����	T��$K�'RJd�DA����\?�@��}M���F��)�;�Aa0��]�[(�`6�M��J3��L�L�j�ܴL�am{���5������*�� ���`V�ʻn� U�/�0�@R���}.��[^�e�A��f��"4I��ҾSI%�y.����.<2�-i��~>��#������# �`���h�H}�`6��{F"㝫�>My�B3_�Bc"��D��J#�NZ�)>&��(�:���Y4T�Ln��1����:NhH%�PP:�5l�db��ܖ��&�G1)w4�hK��iM� q�	ġ�>�8�cQɔ0W��#P�l�Qk�~*9T�|׊`ңb!+��
�6ј����ʷR``�l�}d*1Q��*0��^Y�l� $[I*�ϝx���Gj3�K�����K�=���f'TN�e���%@���¯+�F�0�~<�>�*��${�If"�A0�"�h�l� ��9cS�8C��غ.�}�Y��0�-���{�� Az�XK�q�H�������}��~{��WH)#첏����9~�8I� �S�<���$>0���m�"T��4.�h�{%{A���"8�5�U^>�}��LJ�%-��3�}�"����5��	ܣ�����Vz����q7T����Y� �D4�+���D��@���ώ'�\u��ĉ�%8�7��ܙ�yB�D��^�"�Ї����f���Q�z
)$f@0��2��p��&g*?��D�`�
j=,l�@�h��=yY�q(F^�qE�'9
V�<ܠxhs*��R]�>����7�9��!<��;o����\F����Ss�~A�0&�t�̦^G�v=�f4L���ͤ�e�k6/`������I���"bN�,1oDŭ����,i��)��D�bɉDWZ��HD��N� 0r�2 ~p[�je���v�%����;�>�p��{P"̃.,q�ߟ!>23�Nd�?�v�ݿzK;S�>��mf@|���1�z�F�Z���	�{M��۰�^D����@��_�O���{_�ջ���R���K�e�$K�J�7�ΐH�IR�G��sFs0;9k5�ASeTқM9$��q4�U�����Rjܻ08�Y��Ⱦ"�'��Bs1TQQ5� �����EUU���J�hmʃ�"b�����nT�1y���t��v�����Ȟ���.,M��:�M�%�$#Aԭ�8.A���3*Mp� Ҧ�j�*\�e��ݜ_"| �b<��D)W�x�_�]��BC6�b�