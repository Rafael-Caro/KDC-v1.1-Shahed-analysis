BZh91AY&SY$�gC <߀Rx����������`?zۜ,N�:i�F�$�H$��)�ɔ�iz� ��4 �&�b���hh4z��A� � �`�2��i�B
 d���    � �`�2��H��h@���yM�4������FLh J�>,P &���$�4�'	&��Jx�"�"� BT#	���%B`�F"@�gɶ"������aF�4H�D=�>�M��_,P]��`΂��W��_�d첫(���9)A46�gU�0Vm���IT8m\�-�q�q�j��ZX��P����{�Ŭ�[�p��΂sR4І�]$
��0��$���.���p�^B�a�^���#!�����{���,�7��	��\�"�G�0��,Z�òE԰M�4�cI!`��YD�F1!���
��_,�t��$���/��T'2H�����F���n5M%�4����b�+CS:�_K�]@���0 �@�I_ῂK7Lh`�����5J�d��m�M�NL���bN�d��U���db0R�J˾/!Y�����'a;)����1]�G� ����YB6��W�����{�W���Ϋ�<0:}���[aF(�2�0?df�l�^a+k4�W�����>v2�V�8M��(W����O�sŽ��?�5�\*�������qU���;���B�Aa/I�������dy�Gj>�����ry��
h��R�p�h���7��w�z��i<Go�5ȩ���/�h��5�����#Dɵ�u^�C��SbPR�S�9�;�_�0�-�[깹sN�R
��j���U�đsbs�H�HP*9���j�<��U�N'ŝ2
��q}�tiG���թRI�Y�w��i�\X�L�������R��ciȊR�X$j@-�R���z's��)��쏹��$��]T�W����Eħ�>�$X$q��a�Y#����%V�[V�
��L�XC�T�H���M�b���Ɔ:�_���ģ'˔�5P��'@�z��&oh�li�Y{4�ר��b���t�C�-2X�P��.rxd-�b�&L�q"2 ��PH`�$��k$�1/���d2 �amw:�e�+��	���JSK]/Q���0j�9�B*�,ԅFAJ�����4[9��	3:��}_��M@{��@���1r�Y��t&�8���7a���t����A]��_
��A�~S-�&9Φ�)>��̒'�p���&r���	�t\��1�Y8x44Y�|���%&L��d����(�������22ey)�n���da!r��@E(hW))G z̴Z�m�B&[vfh.>IHt���k��yhRd��6Ս��2U,kHm��`�6+R'5[��}� ���䎠��H����f:��F���J�l*Qo��L�մW^�F��߲O�LB�x �а���2���"�(Hf���