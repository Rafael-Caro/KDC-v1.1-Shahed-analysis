BZh91AY&SYoU  �_�Px����߰����P8�6��Z넡S)�)���T��&&���44 � �A	���f(d =M 4dz� ��&��i��e<�  ���4�	���dɓ#	�i�F& �$�556F�4   4d�|�D �+C�A�/�(��I����,i.v�ңV5˭|�,��GTΘ��=l���t����3�B���_��(A�K�ئ���lЈ�b� �ӄ:F��^Q|u�e~A`��;���CΙ�y!F��J��i�"��۠�@F֤�{�fF�4�4���JX8\ �p�7��m;�m�3Wp�Z�����8n���J;�}���Ṕ�B�a��8a&�-i>R
������/�΄�g59�I�ei:s��N��|׉Y�C�#8���l����%Lj�P���V�}�@����)�S%i��0~ ��6��4��Ԣ�Ť�o�c��(��!�Xz@YPYA�T�B}v��C*z{��ш�|����3)��HtS���<aG%9Ԇ�t�,q3�]K�ߑ��8RE�i���g	ٮ�	4k�D�w�a��,��`1��IE�!�"r#�*v�'Y��WJ��54(e�:l�i#31{ʺXg�j�&i�h\n 3V�`A��\#����!i�w�Q�{01����M��5��m��eqjd9�$��_ŶFYPe�=,ʅN&.+����̀lJ/2�V��z��0!��H�+Fa[���Ӡū �<�Q<? ��h�0�4hR�u	��>���
���j�aŤ�V<#�5S��p���R�S5v9{�Vъ�����ض3P�E��w$S�	�Qp