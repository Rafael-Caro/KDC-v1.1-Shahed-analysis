BZh91AY&SY�Jl  �_�Px����߰����P8��g����	$��	��D����@@��F�OPm@��   	M&Hy5<=FM  4P sFLL LFi�#ɀF	D�	��������d12d ���!A\���F0�l�Ci&���$Y��5V�Z�[p_ ���zH�L�/C�ˬ@�㡶g�$���f�:Ȧ�����'�Ē�Е��ZcSoi�(�x�W�4��7��K����Y����5��RtgS\Մ篊��0-���Jpy�Tw�������cCn�����sm�k�����\�(qǞ#�I(ݭ�y-�f`�(����8�&5�.k�q���ؓC�b�aS��i�i3�j��9�Sk� �r�q*��z��1��;}��Lj#����K���Di~9�g���Z�(O��řW�6�?QoeN+V�Z�.G�	��w��~MBC�Q�i��4 ���97��zL���Ӧ�F��â�~��we�$8S���G6hQ���CM:cq3�eK��"<{�Ĥ���Q��'���*J���QF�-rX2;�����,*b���iJ�S�/�2��V��'͗SW�C����`S�,�b��+��z�o2܋�f!���� ��$�bf������ k��v��ʫ��jhs%w��\�9���Z��̃ a�"N��q<��D,#3]1���%y�E�hݍ�I���F��f;�I��?dݏ<�	9��K ��n��.�G�0j&��C���Md�2��i⠔����)���B2Q�"����.��IRu�wS�ط�XeE��w$S�		t���