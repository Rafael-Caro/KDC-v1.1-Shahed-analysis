BZh91AY&SYp�H  �_�Px����߰����P8�6��ͮ��P4SѦ �ш��h�� h!4������5��h�C@ 	MI�H�bi<��� ���h�A�ɓ&F�L�LQ5OT~�����h�����h4d�%�$B
��1k�DB�������P�cIlj�*�c\�k��d<�}ft����e�5��&w�6�n�B��"��3Y��dN��B " �4""��sf��$���v�^(�
�o�������gIJ=�J�i	�3����kc͡��&'�r����%���ʧ.n���ӹ��4��W����������g����ʆk��FI�	0�k]�G39�ؗS�΋h�S'���s�T��u�����˰��	�*�x��k���otʦ�6%��^ZB�����I3�D�s.^���~����a<T��6�>W�%,|��N��.$A���ґ�CB@�'J�nI�==�xh�h�|��Ws�S��$��OS��3�
4Q�D4Ӧc��^Z���"6�'��-]��[�E:�!*��I�)��72Y=Epe�r� �"�� ӏĞD0�c%u�HL�9�+%���̠6�M�!��3o����*Ƴ	�y5��Z�s�����$�F�L��8I���R�v]6�@�R�b.*��Ps'm�@�]��-6��C u�&I�q�������\��;�5ɧ�v6�"�i*��B�*�g LJ�=?e{p @���P���m�,��B���'�Q+*�5��Ԗ���P��r��X8ba�5�܄�#E.Loz�&PDö4�����$����"�(H8I� 