BZh91AY&SY`r� <߀Rx����������`<]�w���oX{��z1��d%�45=#L� 0��	"F� %Q��2dhɡ�@�A�OPM OPɡ� 	
SM"d�jm44���d4�& �4d40	�10�Bd�O�6)�?*ze?QL)�4� �X@�"Pԃ��
� �B(��K��	5ޮ���_K?mb�m���j�>�}�X�#!��6��m��_J�b�0�F-	�BU�k��\�h�+�v�Τ́��~�s*71)�,��(w�.@��҃��$^�s�B�B!�1�|F���GN������g��n���%[2��A*)P��#4�)礊ؒKe�	���0SjA
�Zg�A	�V�����n@nqAA�����1ǲ0��3XH�a(�
aP1R�)``{�dDJ-v�P[�w!8�Y)��>VD���;e6^��a&�4f�@jga!�*���T��gz�d�+��筳���������אcq��g*L���{���QS%���(�{J0|��]���NJ���gJ�S��b)3�f]cxٙ�4Q�v��/j�g�$)�M�)�/��]��A�3Q�]���?$��_vT��*��\�'V]Q�]2��ݛ^�Ԓ�}�+��=+�^�%BB�y�:z���l�{����O+N�>Y�z7�[U�E�wj���<�:�G��kq�ww�<���?�w����j!� ��Zǧ}H�T1�=�6��<VQ��ja��3Y=���c�^�tD��a-�sġ��	�[x�"�
J�(�_�Y�$֯4�|�����E���:-�lYAMMV��ҙr�5�n�G�ף	�&�w�q<6�0�m4��jN�&�T���8h|�~������"v䬊Cp�/'�mɘ�L��"�� "���{�H��f��T�V�U��L���g���p~��C+P�A���(W ��_}[��I���]n(�D�!J���G-�={�������I��x\�V�V���7LQ�5sE~�CLlhc���>n�u北1����7�C��a4�Z8��<j��9׀r-D�X �&���Q����X�SYō4��Pc�&�2�e��"����D���C4N��Q�22�i� �]��"���*D�2��[̧[�Y��HD����;���Z�%e;��"�]K(�γ�A����\L��H�M@cf�a�ss���	������^�����@���
a��x�ÛwYtܥC���heВ%zp%�4I�`���fG����Fv�[�1X� �+�M:�ʕ�d�NF�I���Uk�Yz-N`)"pzƢp{m0QPP1 ٕ�WObwwz�L��3:���\�����K��+��э�E���4���+�Nd)�[G-�&����;B&���$#aХ�5&Z�3%4fP�k�j�h*�k]WZ3�nq{�t�}Ø��pLE��H�
,Q�