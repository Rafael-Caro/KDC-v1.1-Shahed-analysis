BZh91AY&SY6�n >_�Rx����������`?y��%��͊h���4����5=56���4hd�  =�4��20M0� z C�0L@0	�h�h`ba!"i&SM�i��F�  ѡ��9�#� �&���0F&$	����~��&)�y6T�ML����ʂ�BPv���b�4��%�K�Y&����_���ֆ�m�.�CT��O��i��9�b1��@r1}�]�CBJ�P����������� ܊L���f�c!�[��.��
�uDMV4v8�/��7[f�ݟ�i�!@�D�s�A�|�AT���c�UmF������E�M���AL�d��]xLƉ$�.�!i�}��p�"��ɞ7L(����V�D\@7����1�f�D���a������3.K�0�x�q�#����&QOj�;����2��;�@�dـ�v��y�[���9��j�ū��(�	�i�:O��7}���E�X�D�d�oN���G��Dnm�xRdT8o�w�
*ҸߣR�������L;,I�iE�4J�i��T�^������h{gz�Y5�,��V*�a�Q��ș3� ��B�c��wJ���D0�>Ř�ƕ�/:�K�+|osEBYk�ȁ�OZI���fe�O&H�֍W��}�g�#�Y�VP;<��e�i�n���Vf/��{=���W����<@�`?н�.%�9lH��3դx#�8�6{j �O��8SG�m����q��� ?�|��_�"c����f�5���2&b�Mb� k��G�D�r�����>s�lJ
Rj{�>��C2F<%Ã�����h�׺;�v������z�w���&e,�i�����LٛUim�w(0s�I�CE�)�!��e6��"��i!9	׈KxG��^�Hf���2ISSHԀ����oo3���ug�Hʀ���1�A�����Njݗo��%?t�ܑp��b�Ǒt�Mp��)\)�	�	���.$,BK�E:�	w�$�W締��v8>���ݑFO��X�hbK#�w<�*�ɣ��H%�u�ܽ�4q��W�Ƞb��F�0ar�����-��V�cM03$1Ĉ̀fZ2�C�K��Ip�q<B����-o!Ю���b%C*����S��%6b��vC0.t��ב!>�S�wR�xhL4҈�dlЅ[��nyN��uHJR����ְ��u�q�b����%�4�q����,|����1���n����"y'	A����		�������a������lZ���+�v�vI�-�}��:Y8>��]����~�܎��
��B��@E(h���l��3��ǂ�����[�m��%�hY"�y�������/bƈ�X:L(�25�o��M,21đ�,��]���5�$zG"����v-��ELjmUF��.\�9��Z͠��v�ώ��w� ܏T�U
v�b#?�.�p� *m��