BZh91AY&SY�'Ku <_�Rx����������`<]�<��o0��]��d��S�=zj='�P dbh4�!I�ɦSD 4   h ��MM��244h 2   ��5OM(dѣ�=C@� ��2dɈ��	�����$P�4S��f�O�i���6�S4��6�K�Jf|����B�"��irY'-���_��,���I��k��0�S��r��"��ϣlF4��/��f�2�� pW���#y;��b��b-A�Z�k�VxP��:1�R�����ޝ���ŚN,8
La�lhP��s�X��\"��L#�S��пl�ֱׄw����a��6Ȍ�@�{!q$�Z/M ��w%�Lo	��}]��F1�W����P��=�����62�cD
{��)��v^��v�0ɢ8֢J�H���u@Ԇ\]�SQV�RTb�jG2р�&� `�@B�^��Bb�I��с�ԆJrE��ʳ&�������ᱜ�7m�wdT8u�;{j*�q?&�1yL��v;���iE�cq�[8U(�b*j���=P�!gF[�-��^�*�
HSb�TS_b�1e� R ��2U�O�x���[�fݓ�j-�{����gE�mn�q��
[|@��SD�:,���"�1a�2UO��Lb����fp�6D�V���q85��k�����\��^/���m aO���� ��D��p���DO`�9�!ޏ3eCɈ<�SH)#ⲏ�ÍL2��'�쟴y��H{��j�C;`ж�E���Q�.���ekH�1'�M� wbk���5�U�*�l��-	���7b���$	*�ª���`� ��i�ƛPyk�3U��l��`9zh�0�{��9+"��;��ӕ3�ʙ)��)kx}jL�5/�9�e�&��� ��q�;��g����~��K�P�Y���Pp.ظo������I��d��QP��B�GyT���;4������CBxP	�$�l�o�wŵ��e�i��t9_���yc%ǌn2����0�w!�M3kG6�G�Wۉ�v�ѳ��88A�`\A|L-aR����`�h*���4�YI���@f��\H`�)p��)"�.܉�`�8�F@=�o��835tV�6����[��S��U���QVA��7o��iО����ď�ѭz6lIgY� ӏ���\L���;ڀ�͋A�rj33�Z5�87Q��)s�%āM���@�}'/9tܥCWA.��ZH��� �`lI�`������[��^so��`
x(�J�4�,[m��I����hoَؚ��Y�v^n��P0QtE�N� ��)���� ��U��QUBENpm������|� �� ����E�+���s-	%m��;*
�7<�144ר��9TJ�*HF��K�m&Z�3%4fP�m� ҆�(�
���5֌���/y��7Qځ�2B�8���rE8P��'Ku