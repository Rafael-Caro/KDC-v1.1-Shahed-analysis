BZh91AY&SY+{S  @߀Rx����������`?z۸0���ؠ(��Jy4�4�S&�CC@ښ ��&��7�*i��MF�0�'� 49�#� �&���0F&��5#L�P�=@4 4�`�1 �&	�!��L���&��a'�=	��F�&�h4ѦFLn?t%B�	� ��I-_*���NǷ�n��_�� M+�t�P�I\L��HL�[b+��@yؾ,.h�BN�P�C6�(Rˏ�y��A�e�pK�Mf�ףu+[�o�u��n
�+U�e\[3���z�[�;��b��@���E��@��$�PoB��\ ��B��p��K'�eڃUU�z��2TI�g4��$��U�z�%�v������Ld1���������,�7��L�&>��"As�0��/Gu�d���D8k	Jc���|��1���eF	O/j�3EqpRt���@6�ԍ-˳LRFV�abI7�LU缸�|�/b�-q��S���R_�θ!i�  �أ�"�y;{t�����J	H�y����6VQV��EU\��3GH�x�����'���֬��V�=U���F�4�0��㉓0�����PD��Jg������/���Mƕ2��ӿ빵i=��.����ӟ}�.rq1�h�0w|�Bvݢ�$񐬺O�b}\Y^IB>�G&�/���|W�a{�m�XQs�e_7`3���.���6$H�q���=(���]�w'�KS�}$[�8����K�Z�3>�b&�]h�p2;��ٲEM/����F��0SX1H�8���[�U���G�yM�Au�S�9�;�0�a�[z�|*Sz����w��h������򅖱vL,4�yPc0q!��2 �Y^AsQ,%V�I-�!f�H��A��>��"��y1İ]�I.`���k!��̉%v(�����]�g�q���#��)��cd�	��]��xٽ��P��'���S�<K$x�a��*R��6�Y�a��^"��]�E���r~;o��i�c:�_#���s'��,w���B�74r4i�l�Z����xrq��� �23.���F���Z�*-$ƚ`dHc�� �se�C�%�Sa$��� ��0s1���k����VY\�_@L��2R�[.�GɎ%6`��fC/,p�զ�1B|&.F�E���:iDK�>ۂ��ӗ�h�į�ER��CVYl44�&����~F�m.�]A�It�W����S�f(=�e��s���O�5�$��%�9�gL$H&��Y����F��u�`��Bóvʶ*��ەY���G[:ߪ��Jm[�F'}��da!t��"����C�=�Yڸml��#$�6-�\Iy�*�D���4���Z�T��3����&��j�ҿ	����_&���:�F�"ۋ�u+����hkTF�K����o+V�YR��0�g��$��uD ؏�Q
u��#/�]��B@��L�