BZh91AY&SY�?�) /_�Rx����������`?sw;ls�'N��C%2hh6��yL�Q���i�4A$I��ji�M��  444	I�4�@ё��     �&L��L �0L�0�2d�b`ɂd ф``$F��cB�MG�i�i�b=A��=M��}��	A�O�	� ��I-/�"2����|_şF��m��|ړ�O����D����؊_�H�/4U�Z�@"@/�J��7<��{/A�S
���z�g��4+v�&G$��P�.ߓ�$�g�����Q�)m/)wT�*.0�H����[J4X��_ȃI��lwI���RIu��]-���7�zDa �d�z����y�<�)�CH��=�҆�J��E�H�4��љ�-�
P��J�T�(1��R��pI��	3`0P���P'�;RCQؤ�kC?4�A�f5aR��+����v���f��6�l�d)F-�[H�֒��m�HV ʈ��q�E]�VA�ZVO	VΊ+;U�C
B�N��)Y�We:��<&�Ld�0Y�ś(o��f2��]�l�ߚ��)=/߾|����>�UI���^ƌ��Q��a���:'����ъf<\Z��h���c�I �$B7�etX6�s@���]۔(�L!�|��N��s�i�0�Z�2S��v����D�M�$uђ;�5T2�� �OL!MK4�1U2f��k�����a|#�Dǲ#�km��P�t�^4L��Mbb�5��#�"p�������܄E���r\lZAf��^�^�r�Ω~!I�6�p*ȣ*0$�L�8�qE�i�ƛP:c��sR�O{8�(o��
dʎ���Y���GIyn�4�e�ZT�L�U������!�ؿ�bA(��	�豤�6��冉����E�P[��1�A��.V`�����"�S�$T$o��Q�U#Ӷ����KXC��v�	q��;)����2AL�����CK�}���,d�p�#5�"W��S��jf��憐K�W�)�{ h��.�!��X8��2#F
�F�z"͐UIk4��I2$K ��2�!�H��C9$��� ��0s1������ �@�*�D��pL��2R�Y�G�Jl��QVC.*l��F�/B{&-��?>~eϫRKEm�0Ç���W)�ȑ��l԰�<�E�����j�bn�iy��K�5�wP��[���1Z�:��nd�;Ӏ���I3��@0Rs�C��S��b\����d
YQJ,�sI�'�g9bNJ���L���pSj�w^l���UE�.�t�񉒒�����c�gm����1L�.�η�xbM"Iv� k��x�Vd̃&Ս�B�V.kWܑ@�*\��*��KKM�A�M}�A#J�]eI��t)�F�����h(X��(�
�nkv+�|��'���:��zI!a?�c�rE8P��?�)