BZh91AY&SY
w�o ;_�Rx����������`?zۻ��l��s�uB+�I"42O@��4��OP6P�A�&�M�PQ���  h@    a�~�H٪zL���M�!� ��04�"d�OH=M  � h��2b10d�2 h�00	&�MLMBz�SOSM�mM OQ�4�����(9 ��b�D��KkK�,�w�i��Q��/���	��l�@K�D��D�i��lE�{d�/4Y�R�`��gDm���ͬ�m����261[�|�����䶜�4<�\�0N�B+Kv��6lf]��z`�����`J�Z
�'H:�Zmy�ӣڷh��2�� w�,G=	�H��[\�Kz���~��g�MIX�q[7MP�g迷��"*
��^R�A���Hy0Û�0 GS��ct�UvsD�Ԩ�&.<yJ0\j��nsA�Kw�V�+�((�u�Ef��E�Br�,*�3��@�[��#�f�Jd��L�]S�z���}.uun�@� -�a;@&4|4{K1��\7��� ��*�oY��pRb�6xcV5hxܦ��!�ѐ�]����ɬ0g}�X���J��	]Z�;����11�+s��%Ǘim�HC�8��|�G'.���!:�r�	bV�&t�,p�Iێ�a2t�&�ᛯ���m��me�)�8�h1�{)*���`K.K��娛׻:����n��x-����=@|`<�Aa/�����;���vg�|{�ڈ;���
��-'�͌����G�鯬z�i(>1��l��n�a��C
�)��<�(Q��cǥ7���X�$ά�������ńa��|�R�,���#�_J��e��C0nFm�;
X�Ş@���)�Ƅ^6Z	M+��
�����'^��AGi�^��5�,hP�Z�R����R�{٨���U6���_��&wiW��T�\A]G���Hp]�뻂�����%I�m:\��'�����d�?D��,y�w0�]�|9ֈ���.$s����4eӈ��w��������\�y�Ӊ��$�r�j�	�����@�4/m�˨F�t"�\��2�2�X��hy�.��ʫl�����H�@3,�p���J��JE\a	�d2 ��nuu����Nr
����[.�G�MK'��19A�>���	�H(�4ĕ#�͍sa�J�!d��O���E� 8�72p�1��"�븼�L���a�jd���2KH�l=|�7�����t��җ�:�u���"�'	A��1��	p�u���Th�ij�,&T&����$Nzg%A�akcHw�m�(ݯ�#��r�1Yȼ�y(��5U*Mc�{Y�lX�w��9q����AbEIіL�-�]ay�3�C�&F�G5L�a��$�����N,M�5�u�����X����7�0A��UK˖��/8��*��,p��l��Ƨ9��pq �$�zDW�rE8P�
w�o