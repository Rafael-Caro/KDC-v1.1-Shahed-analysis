BZh91AY&SY�(�  �_�Px����߰����P8��s��Z�	$�H�z"z�D�OSL� @@�h4
dz44 ��  $DMRz���7��z4OP �=@hѓ �`A��2`�HSU=�e�2LQ��5�1M4f�|"D �+v�A�/�(��I����.i-�U�V�k��|�>L��#�3�n|S-qXui����;s$��w��
0�!^��v# ;��I,&Y9�MTӴ��)��<4�잁b����'-�t8q�m)G��Z����Q1��"K�:�8�mP�3�'��U�Abf
���Z�w�� fZ�e���8���I(�~�5p�f�`���3$݌�� �]��b�A��>dw�D�7��f����Կ��c�'+����ϼ���ѣ?�%�5��XwC�h��D,[d3q�5ɭ*P��_
�����2�$�2�����h)c�����1EI�F���H�!�B���y�&�:5��C�Rْjz�Q����F֟��Y
8h��i���έU.W��r�H�(�����T�"�'�����3ʊ����<d$V(zH�B3�#NDQ%{~��LN������,�?n��Gk������3�V���VfweI��&"�ц�dë�A�2On&yJ��|ٲ�U-w"�փ�2�dE/3&}d�l{��q6ԬV�s�������ch�|j�}[r�b0��=jT,c0�q��(?��f|�&L	�
�"���8�1��1�EA�/P0��G��C	���YL8k�f! �*���roW���l��q��:�6$�g�3
�+m�I�.�p� �Q�