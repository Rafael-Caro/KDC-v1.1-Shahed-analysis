BZh91AY&SY�m /߀Rx����������`7|�4�u���4h���T{T�'�#)�?Rm d4шa���$��)4����@44��b�LFCC �#҄��?J=Cڣ�@�=4 M s F	�0M`�L$D�ơO�h��i�4i 2l�� {��
�,'$ ��A-Y>z�����w���0�c�l4�>��K�C��D�i��lE����/��4,\��÷��V��_?�~�}���P-fi�MT�\�l��߆�K�a��Tc�<��zq�s��k��~ft$H5�ֺ@g�j_�����������X���p�d���<���tQ'��HtܺՒI-�������f�r&����F������FA�`��$$H��X64�����-C�WBU���G����[��Y�:[:%a�2���_-�[n�h=)�8�Q����)oHl��f�cyy�_%r��m�S"*C��?���/��Y�B�H� �lQ�qy;�t��9t�
��6�[	r���l���%�u���R"q��Y�x�dе�C�k�p�j���j
�Uj�J���^mMO�!1��`�e��k.���nZ9l��䶨�3�G�VZd��c�C�.Ȱ�Y�S,#��b5���������$��*��Ԯ����$G-�˗g�nlWup*����[�4[��x���\@�lH��.��Lz��7��ڈ<�[8TG�k������|����X���%���m�d�6�\��(b�Qb� ��▖(�	��v��u4Q�Au�T�Jq<4�ߒ1�;����ts�H��[0�4�8$�^���K>)utذ��cM��4EYf��N,鐰j�'�[N�{yI:���!��2+͞��[ʘ�Լ ����!�ؿ�`A(���꩜���c�q��~>�&WPWA�cd��8���[��@j��Ӻ�.Q�IƂ���#����%�ƅ���*xOIBTE$7�L�G8��tW��-�bp���v7>'��ّs)��8��1'#�x�f��ph�mi�`�����F�����Y"0�H��B�����Y2
)- �&�	�H�@3-,�H`�%uX�JE\_	�:�d�B�� �Y�+�7��!)3D�]z��M�P��
Ah����B�AI�"�5!�����i�;p��}3�Ն�Xq'��ٽf#V����k3�!���x��K�4��A������4���4n�1��,l��|�"�'	A��3�� )9ϙ��_�F�,po�d�,A���c*ت��nf�<��K]T�+��G���Ks��"�+v�k'�LT���6�i:�'ww��2����|��$�$��4�i<2)2f!�h��|UKQ��x\��+R������y��}]��A&�&
�v-��
���kUF��ˇ�fZ͠�V���g�~�|�0�6#���I
���F�w$S�	 O���