BZh91AY&SY�p��  �_�Px����߰����P8��g��G0�Jz5A�����Q�h �	(F�	��z@4 �   	�H�44M=&� F�P�4d���`F�b0L�`��)�覞=M�   4cD�	����~(�#(_�Q���a��$Y��5V�Z�Z�/�g�d=�>�<��|L��q�����٣<���`Q��)��)]���|�T��i�,�)�4'R3����K o����������6��ZBn�Ǯw�'=��%X�4�I��ЖO=��������R��=CN��d��<E���\�(q��#�I(ݭ�x�����.��M�I�`��r4���.��!���iN�(����f�.x�����J�ޜ����;���T�%{���M��G�q���9�1��9�򉶸՝�s������Mj�%��,|��;?��>�e>�D4��
��o��eOW5:h�j�|�׫�4)��Hl��߻��F� s�t�,�g������:��Ȥ Ә-�M(��bU�1��u����7���--b+T/I5w'��tɨ��g	R�T�غ	�UC_�d�F�n�K�,�la�eN����J[qRV��>���(@B#!��DTQ���f'�#<�D�|��[�K�d^U]t��Κ��hݴaq�l�T�Os���Hd؋���P�Ɗ��!iJ�$K�Q/�19۟躨 �D����`��,3D]vNyEȟ�G�9��6�
-n9�i`���E�G�Jڃ�e8�E�ı������1�Ωf]�{�#8@�2.���"�(HZ8EQ�