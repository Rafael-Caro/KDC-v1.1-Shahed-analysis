BZh91AY&SY���� _�Px����߰����P8�7L�j�Q �ѧ�b@mF&�   ځ�L�H�j6� ��4�b	�������Dbd  �h�A�ɓ&F�L�LI�����2cS#@4 � @�!AZ5���a~�F��M���(H�����J�X����2��z����7<��[a\}Y�wf�7�I!ye"��3#j䭜ȶp�KC�J�Vg���yͽ�`�0ϳ�FxX,U��g�/7oK5t����+h�r����f���+����/�N}�֩� d��	���ߎ]�m�t�,m;m�3��t���t��ZIF��xV��W�pζ�&�dư�%�dV��.�g#c�5��7y��Bi��.������Lh�� ��V���`����`r���s�p�Ψ/�H0�wg���D�����K?pZ��A��n"0З7�RM�P�>Y����)D!�b���Ă�F�JP�]�%ES�ݧ��F��ǝ��M�<z"Izz]��(Q���CM:c8���`[[�G>�����a֭6���R��ux�cN��O�0�k��)idrh&��k��ND��Vj�Đ����I�
�W^T��*.��8���S�Y�*�q�s��m�����Eǎ�i��`�A�d��L�*'e�kdi�]�qUm�mM+�q3|\g���Hr�%��_����ΐ58�2��M��SS��ecщA
��Vo%:�t����  ")]B��0Y�A離�`A�`��"��sfK�3�ݜ���%c�Px�@+)�{ENER��~��m*X�z������ �B-���"�(HK���