BZh91AY&SY`�^ /_�Rx����������`?y����s�:�:!��4�0���h�� �d���
f@� �@� �� �����CL�� ���  �S$	OJz�=G�CCM �8ɓ&# &L �# C �"h�4�S�O)�MM~���i���i�LL,?\%R
��(HAQ�Y���ҷ���\����D$�U*%�WH(f"	�	"���9TPd�Qhh��uL�	�o�`�kPiV�Z�S#9�	�#��	e ��>I��$�nWa�H4����b���� ���^𔩵���`Jpʬ_�u��\fٲ�"�\/�.�<�K/���s�(袒j��x��6��"@� @��6���AlA����D���"&y�8z�TFV�
(1.Td7"�����&%�b͙
KlɌ�ť��f�4�WLV֯QJ�C4$��9Q3z��%�,q������:^ov�5��6��hlBM$�GBH������q�]�/W(el�xn߂�JK�T�Jm�Ã��N�C��4"���qZX,���b��iPa|]%٭�u� "	ҦJ�J�/-��t��W'B�33;����6�7lC9���Kl���vw�ˉ��>TŇ�����t�9�_tbG�2�b�9�����kh�,�LA������q$6��<ky6�y�;��@{��D�=��!"G�Z�&1ޏ�������V�
h����r��_!��� yi�B�GD���#��m�$Zgt4.�h�{5{����pH���V���W#d��s�[c[�9�(�$Q}��ZpA���v�X8��Z,�7b��D�ZڱN�ȉ.�(HP�0P���Q4tԍr9�%��`��$v�$
9����{�2&[�w�$�;�jP�l_&j$�����Fd̭�v���s���T�,����cd�	��.�4V�{�5ȡ)�[�*8�S��*���zKV���{�G�|&B+"�l�n�P�	�`�Z��v�_��������W�X^K�u<�f4L���ͤ�U��l^`7w�H�/��F%�0�Q����X-mUrcM05L��@3Y`���Iv�l$�1a»�PMh`{\l�ۅ�Ub%tA2��Jil���8��{PD���U��DAJ�b���Il�l�rL�=$�N_3�殳 =D���ٹh#^�[��	�=�%��m/]a�Ir �qI/]���Py�a�oY}�i���heВ'�p�pnI��"A5H?���]��`up�kX�� �U�X�Ni2d�6xKrTp=06̍L���U�Ձ��X��UE�)�Ya�����r�Սm�j��Y	7R��tC7� Hy8n`�Z�J�z`M-C�Ⱥ�y��c���4����G:����KA�M}D�Б�H���h;Ko���r̕�ib߾KMmmU.k���{n�O�\B�P2��[t%�.�p� ��"�