BZh91AY&SYj�_� _�Px����߰����P9������	$��Lbh	���T�6@�#	�	Dji���   �  �ji�ړGꟐ��z�� ���4d���`F�b0L�`�%=L)���D�    4]D�!��~��"�_�Q���a���*�]�iX�Z��s��D}�l��H�`�����UL*hL�Y)�R��%��dLp�>�J�~G���6�>w�L0�e��Ez��o�K����3=�(���+h�r�mL��M�N��n���uU%5�qVaB�i��վ�M��WN����1�к�N�8�#��Q�?6��1K�陆�.e�}��[�diX��v�d�%��Y��:�-����W'���<�W�a^���O�x�g�y��:k��+�o�}۽C�H��sj�sȬ��aQ�͓J����J4�jSgmj�ʘ�w�X�)���tVj�z���	97��B4�g���/}��C��/�"��h^vXB����4ӥ�W;v�T4Y��y�D�4�㌦���r� �S|K�TgND��s�� Ճ,�� b��]���Ր���Ul�/�ʂK<��^+1Pи�3��k$"iib�!�7X%�kH��i���*�@r�ȜD�F��ɇX\n@�Q�M%�Dr,$ت�-z%�BC�1a�2,�!C�i[�D���� ���%U�g3h���9�� _8�"s`�F0lb1�%���F�˼05I���6vm--В�RB	ט��`�7!���E�Kt�#���6�v��2SQP��� ������@��W�*tU�:�Y��#�mU2�@�HG�]��BA�9|