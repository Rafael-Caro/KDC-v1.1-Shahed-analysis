BZh91AY&SYs7�Y <߀Rx����������`?zۜ�M֣��eѐ�	�Sj��6���4dhCL�@���F�0D��i�h2l��@���b�LFCC �#҄MS�C�ڛD�SA��&�� s F	�0M`�L$D�4@L)�)���113)�CMi�x����s
$ ��J[Z_
����_��n��_��6 �VP�%��Ԓ��#1��m3�m�����b�X`�v���@�p�Y
}�2	�n&���#ʂ�m+�E�,�;<�M�W�Z�1ڴ׳�������ʚ���Vx��v1�s�I��AE\F�ܲ�{��B�V�J�J�0����Hs�v9A$���/�%ǆ�_z��됍1��ۧ�ǴFav���D4�~A�-.�hã���P��T���5>����0�D��5��g�WSp�]	�&b2x�w4�Ԃ�����XA:��r�����p��,m����V�_�Ĵ�B�D � /#b���ӟ����N�҂F�+]/*����YEI�Al]�/ �K�FP���^^PًO]1� f����PUb�VUg���jx� s�I�٦��7�(n1���ʿ�^vW��Z�6�S��k�K奖�Q���F��{zL�q0I���>�! '��������e�?���b���36�/��Yb���[�4[��{ ��{��Aq/9�C`2C΁p9���߈W�����\�ڴ�9ni����^���sIA��=��l���`+��1��LLR|^I�Ѯ���8��4Q�A�T�Jr;��c�2�;�6��ts�H{v�\7n�]7��_H�'������ZT�m@4�1e��E93�B��<߁m:����;5�%!������3V��ej]�J\��%�T�l_&h%,2AUD���F�z7	������)3���;$ �⼢�Ê�=���J�OM:ܢ�'*
�e�;y���9[�l8X3\1@&}�����l�)��/o��7m�PB�1��ϑ�����`�uuNF�����Z���9ZA=W]�����i�rq��A�ɤ�.1��.��]Um�4�A#Ig��	D��	H��a;AA��?[�D�2�N0tJFL�-�b���Fd��9�H*��B� �L�M���Nn��N��.|���1�`:Ǜ\�p��X��y�A�\N\��FM�m/]a����-���m�H���!�wY�])cg��`k�I�8JPoI�L��A���яm^H��U@P�8�^��c*ت���Vl���Պ�U2��Qṯ��ޘ����.K�$���QA=<�烳'H��ffi�NZ��9��-�	K����0�H�`Qю�7��E�@�.Kd<�)nt-��9�5�v����\��#�l��T��Z�6�0\8@q�ĵ�Au\Z����v�� �A�9�:�!]��!���"�(H9����