BZh91AY&SY\�� _�Px����߰����P8��o]1��4�b5==�j#i��&���M
{U?Q���yPi���0 �� H�)���<�CQ� �z�h9�&& &#4���d�#�j����O��Ʀ��4   2�=bD �+~&�"�_�M���a���*�\�Q�F��&��5�YKdpz�FZ�r�霸im��t�⹢�ټ�ޮNt�!@D��dTA����1���01�e�J���o��'����f�s}�,�nO��8�	˷�J�WLOr�C��/&c���
�L��R霚�WNͶ���t]���B�:";��6��yV*��ܙ�h��/�} �g�q,JZR\�'m"���A�i��wv�����[�nܻ�#	�ݕG��ctz�Q�9nI1$���i�T��@SDy+��PG�^F��V4����1��2$�Vğ�������)v� ��f�^,(, ƪ�P�����.��s��yT�5r�+#C@��l[)>�\�9mCM9�q)n�B�j]�NRW�)��0]n$\�A8��2��Q�)������(��[�.`�?Q\;Jc�J�J%�?�t��e�PR_�mL��m�Z�@��ƥ�K��	t�c�6���iq�f�2��_"0d-���2G��	%4�Vl��K}Q�����2l<f���l����h��I҈��on�r3L^3\���OM��b!qZ8b�A/D�0NL���q�x�@L�Ekpe�ȖY�F!fm����q�a&X�uk
����	��3�^8bq��9
$!��'l�*���Yn��cb�f�.̋�ܑN$�%�@