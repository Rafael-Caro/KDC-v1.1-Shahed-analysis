BZh91AY&SY�w  _�Px����߰����P8�k�l͋	$M2$�hhL��lMF�SjOS@P5S#z��@h4� �  �`	OR����ɔ=C� @� 4d���`F�b0L�`�$�<���j�OSA�@  d�zĈA@W-}�"пl�Ci&���$U��5F��]/�u���>�����=���n���Cl�I���&���2)Һ�@9�
��U��v�駁�섕#�]|w��Y`���$�85<��Ĝ��.M7'�hZ����YLJo��B��=U��Fg�0,�c/�x)i����Y��w�� f��Ĺ_�
r��r&�>�%0`��M��FFL�i�&Ui.h�&/pw|g�F8h�{�{	�U^3��<l����!U�%���4�:ĥZ�\	��'d�!帨ݾ���(�eSS�b���G��RN;�;��_݁��/�We�D���^�(h���,Iɿr�S(;&�3�o�JZo���9��\�ֿ�5c
5���4ӝ��%-�hT.�Ӹ�����S����q����5JFp�\8QKU�0�k��+Hh��=xT�X>t�B	_׀�lT��tV"�5�*�Ls�7���xŘe���oԸ���+S����e��ĄZDb4�\�	��2G��2Ji��\�Y�f����w1&C�lPB�A�v�W�:)U�.s���Ty#mE�c4�=͒�2e�g��7�RB�f�B������H���g����0�k�őp��/D��)2��F�|��c�&k�D���Z@"���2�9��NX�%6��th�1S�.����l���.�p� 1��@