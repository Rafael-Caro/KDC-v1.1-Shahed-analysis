BZh91AY&SYcn�	 :_�Rx����������`?z�wn�\�70�kT:0�D5<�#I�)�T�4ަ��4��hd'�4�d@�Sj� �@  q�&LF& L�&@F �)�
dS�&�242  �4�L�1�2`� 4a�hF���
��O)�z�О�M 2bcA����H,RHAa��4�� 7�u��Ks�t~�d�H������+�
b1�-�c�<�_�
4Y�I����o4���j������b���'�g�����m��f�T8Q���ɜ�돁$mn�/�ے�C^�4��X�~z�G��U�Le�
�2ϳ�ʻ�Lh� � M1h}Ap�1������o:�r�vt�gɉJn���"+`a�l�����l���"��m"��0��//�ydRw�(j(nE'���l�ljm�%�A�h�U�E�ṅ4�1.�VP�^E��)�-&��Rn\�NcmV-A�y�k��:_Gǯ0�&ѱ�JC�m�ϡ&I@�����É��˪F,��L���7ܧ%Kƅ�h�Å,1�%�&�iF�N	�t�Bū�g��X���J�e|.�в���0EL�d��\t?�M
���eW)p�Ngu��=~�Έ�2�2�ڂGEp��w-.�:qR�k<r��~�_{,�b+��:MFR]Q%�w5E4݌z�|$=]:TבKVqX;�Ê���u�����p�H��-棿)x��m�g�Q�=���SG�i��i��o��_H��]L|%/-�k��e�
�/�h��5�^�)��@��E\��P��immn���(�$Qs.ذ�R��q�kA�~��w���K�Tq��n��a�(P��(`�_S�0�i��8d0��^��G�/�w��g��cBeٯ!.����Z�I3Z��Q	SSH�H1��iw��&�6N���Pc@jEuK $@o]���w7�A�"~�8E�s�<K$wq�Ἑ�i�l���r�7ÈnTM��q���/)[���Ӏ��:_3���ģ'��P��NC��C2�f�fƐGU��3Z� ѷ��9�I���w0dR�,1��m�V�cM051�	j$�&PH`�!v�l�Q��,1�	�k��qm�s,���G �$�dD��KԽ�r��L�DXs�4���P�E�w�R=��{v��Z�L7�|?�ٚ� ���ͫx��j�Z[S�,��I�#2\�l
�%�8�b���̅#��]>C
���_a>�ӡ$O�JG�6�Ω$@MVGݡ��K��eN\s3Y�@˕�M9�ɓ�YD�*�~'L�je�Jm[�,N���da��H%J*�Pf8�Ք�⪪�(m�")��p�!��Z�f+!*D�Oc8�`bl��*^J�L0 �,~�pbh>)���� �P[qbb7��� �T��ETl.(�n�o��]sh,�{\��g�~�|G�{���
�tHF/���)�v H