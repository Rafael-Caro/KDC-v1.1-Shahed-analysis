BZh91AY&SY�
� _�Px����߰����P8�0^��+���5'��MOS��jz��I��OSM@�OI6��j<��   �  "D�b���S��4����=L�1=F�P sbh0�2d��`�i���!�J
�����D��jh�4    �l��$B
�V�����~�6��M��P�F��SJ���U����}%,ѹ��et kF�'-�6��/�XSz,��,8�yK��tPp�FNI*��sgঝ����a���۪Y�r���I������stՠ�@$�r{Z _n\�Z��*��$lBj�T�TRȱQ^��g�ҷ��tm�@̺Mek��Z�P�v��3�6��<��*E�ܙ�h��7]"��oh24�I�.�<ޤ��F��պ;z���?6v�p��:wM閨��Ԙ�Q�5����_?�g���;�~�KN"�&5�,��ү����'�'�9�b���ak�[��b�iގ���h�CDAZNM�:R��բ7��qF:�IK߅?5Nx���kJ�c�f�,P�NwEJY��P+��Q�A+��է/Y^\�ƜL�VD�i
}�>����	0�r���-*a��_��E���:��d���eׁ7<��h�X� ��,
�W�%,�ƕ+0O(1%� !0�i��
�2X�JT� ��5Bǒ�(��8!�	�A,�"�Κ��4
m�"qP��4�'����0<��c2�;-SQUp[D,)C&���TK��Į~��-� �9��{+U��g^E�ߛ<��� �sE�p�f룀h�!@�q���\0��$�N�OL�qD���te{_ ����@������H�
aZ �