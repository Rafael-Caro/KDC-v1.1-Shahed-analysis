BZh91AY&SY�q�� ;_�Rx����������`?y�G=��Xy�=�u�	D
0��������P��h �� h4%Oz�jdҁ��� h=@� e4��h=OP4��    BD�i�@���44 �CM s F	�0M`�L$H�4M5=&	<���&��&��d2ba`���(9�T�1@��B
�D�ͥ�Y&����ߑ�3�֍&�]�v��ޟ8,�1�r��c_ր�b�0�F�	�BU��5,�����ㅺ\�����V��5��a�'����I5���ׅ'G���3١���E�l���с�U`�SpW2���v?��
Y����Pk�Xi���%D�+��<0�I-��X]�7%�o&�R`{�_��b1���|}�u�*�7�w�A)�y�	���oP�ȶ�C�_@���5RP�h����)�J��`٭dM2�ͨ>����fR��p��"�#���*��E
g ��^��u�˺���E���o ������"7��:�dT8v���k\Oϰ�f/)��p�SǇw�(�Lg���z���xF0(�Ȇ��[":B�T�Z@�jڳ�ي�TjѥA�	S�^&N� ŐBdF8�&_�U2��Riw����C��"�tz�|��,���H��l���69aҗѯp�ǧ_�8�l�h��@��X�M�1.|�ac�aw�Պ��2�����Qk �o�����.��D6$H�a���=h���|�v��[���YK��r��_a�&��u��<��R&=���rH���
m.�h�{5{����p$3�t�y��73���!���x�k"�en�Q̚u,�ctA4h�(l,�	Ɍ�I�$R%@�HPĻi�ƛPwؙ3U����A�ӆ��(�n$td�$
;
o�ʙ�YB�D�t��$����Z�!�������SH̀��y��~Q3�a�����#�)��A�j��ͪ��od�%>��"�#��:��8Xq�V^JS�i��2L.mar!Zj��b�p�O��r�4�Ɔ;NW���݁c'ǌ�2���0�z��h�����H%ƫ�IȽ 4k�.!�`^!��K.aR����ZZ
�,�ƚ`h$�%��f��!�H����RE�\!�O�a�22�m� ��a�+����X�Pʫ%�|��c��/j��!�7o��a!=�g����iDJ"�����7,S��4�T`��JT!6��ft��ӆ�_��6��.pŤ��[����Ӽ�Pz�����_G9�rx��Z�D�N���gH�MRnG��]��`so�iX�� �����=�x�T�	�ͬZ�BzEڮ�l����B�7���,1TRR4�@�et�4����34,A��
H��_s��gKD���!�͛���W��5P�&���H�,>�nbh?	��G@H�R+��1Gim�6.A���3-,[6@m��[kh*�s\��3�vr{�9�r#��Q
v�o��rE8P��q��