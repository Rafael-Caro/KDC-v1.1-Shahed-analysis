BZh91AY&SY_�V <߀Rx����������`?z�G��s��� �����M4� ���  ����z��i�@�  ����� 4    JjRz&Lhd� �3I� � �`�2��H�&�����ѩ蚏�'���4i�j2���!(;\�ؠ@M!�"Ini~��%R���
sL�fI!���SBA��	�2�i��"�}d���aF���9 ��k�r �fq�〈H6vNFb"9��_u��W84��&��<�������7p�������J	����P�2�V)�w�g֭�L}n���i����p�*��On��RIq^[��ג\�g���5�{m���0c�f�����# �`��o�$��Z�F�0��0��0<�0�����%�΋�8v��ȉ:u����a�8o�a�m��V�f�Fq�Č+:�aZ+����q�T��գAG<u���$����	h�*�}����$"C�!'$�H�J\&���/h�\�HRY�a55�Dz''(��t�E�	������Y8(�=kz�Y5lY��V*�a�Q�H�I�+` űB�$�}I��u#���10];��]�6�<W�;�,&�AxDMbڲKq��s�LX~]7y赀�mH2̗(�CY���TdN�#��pa��+F���y��Ӈ1.�d��h���G�	=B�l=ǵc}�O�=��V�
h�ֲ�1�g��3��0M~�_(�1��sm�l��������SX�H��g�!��Cυ3}E��,&`�dE�د"��{��>��C�$nU����3T(�\$���1P��PZ(�i���N�"���N'ѝ��d�E��D��U	�"����i��sRe�^�$�PG��/r�3j���T�T�7~ؚ���������~�FT������+�.�qV�v�@i"���>�$\$t��q�]#Ü<N����k�g��Aߠ�����/�)�<�ݏ��O�~:�ccC�������d�{e��Idv�Ω�:�A.ۯ~������tq��!�H̦.\b5<=��V�1��	&D�l �l����Iw��I"b(a	�9��d��� �Y�TD���&BR)M-��G���1j�!�9s������)��÷�D����y7�In�s�q���]�5�H��7�"4ٳi��XMq:u��q���wm%�Am�d�������?1���Ʈs���O�5�I�8JPoI��� ��-O��0��2;9�h�\��&QEA(@��I)�I�д.@k��	_�fG/ʊ�tc!v��"�3URR4����C""$����L�P+���A�X�W])�ر�f�3���&F��ULia��$�����&&��&���֤_�rb8�ű����ƪ��X�����%�����f8��O�tB���|ʡNޜDl���H�
�#j�