BZh91AY&SY۷� _�Px����߰����P8бm��v�(�OSFLD�P�  э@ȓM��O)�i�Ph�h�h "@��5OP�S�x��4�=@ ��� 0&&�	�&L�&	�����jaL��d    �i�!X0k�4���m����P�V��5F��[t��a��#�)j�O���\�q��b�:�H�\W<]��.9�ۋԩ]�&T�I&�US��\�1�m����z����I����3_s{zK&���֛Br��S6]h�t�gJ�j��~yȪI�f~��4lǼ�1��m�@���ye���(q�|F�țt�<��!��n�h����} �^�l$2	��,%��s]?(p�F��Q[�)����@���@I<[_n[�#<u��j�s��Z!"����Suٳ�PTY�R�����No ����bDa�#�])66�J���0l��B
���j���TJ��f&B��t�$@F'�.-m%��W�&dk�Q�h������l�P�.ʎ�bW��p��N��64�$��m�B�)��ޡF��,�� b���Tëy2!��a�m�H��2�]/�]*��tD5b�ȥ׊��PI��� �a��ZNf	B� 1~tP"##9�Drp��h3���IM:䕛 kE�U
+Y�i�g��}-A�v� ma��=%J*W1�d��!�8�!�〙�Ze�����^C{���&�)#M�����8p��A�_P��	~�+���l.�$/r��Q�MR�h�i���	��Ux�cy��I�(Yk.�A�)Ֆ��l\��ّo���)��ݾ�