BZh91AY&SYN��� _�Px����߰����P8И�lWvI�Q���i�16�C@@���`�jM?TyCOP��hь� ��	=6	�mMH �z�F��2b`b0#L1&L0JHj       螑"T
�ů�Da��46�l>߱BEm%�j��MV��K��d=}�uF���2�����Iߝ�f�$��|u�ˌ��랺��@0@dDR��:R�hǍ�$

]��t��`��wB')nM������*�	i�}m%{,���x)����&��s����WeW�ǫ R5K^���V6�����i�X��oI
o��I(�_�j��J��f�h��7�&@����9A��򹿁Μ9.���.nq���;�Y�X��N���eG]�}�,8�&%��`o�B� YD���jC��F_�^egxkp~"@�cIŊ�hR�Dh&c;����c)�G0�j�g����J��}H�#O:8�6���D1�Qnl�" ޏKBxь(�Du���0��L�rTVUu���ң��5i�Oi7� �xȸ��v�'���Q�
|�iL(5���hS�0���G��8��(�k��)�
�h^e�u6�DMi�V'�e���Y������ևj��2X�DbB0�1d-P� �2On2��ٱ��T�~�ZT����%w�&n�N=}@>,��I(=W�V]pwrB�h f�bh�K���ӆX���ejX�ųpbpI���5紴�BK�I'V���V�d':�Q� ���(&,��a-a'S�mƐѺ� �d�p?%���
�0���C	�kSF*��η�cb�f�.ȋ?��H�
	��W�