BZh91AY&SYW�� _�Px����߰����P9��h���넒L�y4�4ɚ����������dځ�dҞS4�Q�  4 �&���D�P G� 9�&& &#4���d�#����S�O	�����  2 3M=bD �+��A|/�&��I���
*�\�Q�F��&��5�$}%,����0�,~6*j���Q@�D:l����*�(#k�"ps�
9$�8�q�ETQ�ӦT4�����\�xB$����c���|�	4ܟCKl3&6ɒ�%�8��h��db�1:C�u4xCN�����o,_���B�w�sNDۧ����r��-�3��/�k*n34�E���4���Y=���y�O��w�
�o�1����u���^m$���)�������\)0�b�}]T��ƞ`�/B����&%�8Ԩ�7Z�L�Yc����1�C��`�~�h��+Iɽc��whK�G!Պ*7`Rg�t�����c!F��r؆�s�*�R۶�B�]�mį' 5D�m��N1)Ы:Xg
e��	,�"�X2�&W#�D�X�5d��"K�%*�9R�3�V����jd�ޔ�IX�nA�	��^&e�Աq���{h�E�#�B��4�H��a$��m���5��wj�J+,b�T�f#��Dӻp�f �h�2JR���_��a��0E�r9��^>8�QH�וE0�%�IC����jD�"HI�|6�*��w�!z��$�!	�)5�>��F�`���L8b��� �K���9H����L�P%]�����`�VY��l\����g�]��BA_/dx