BZh91AY&SYĝ� _�Px����߰����P8����0�H2(��
z�SM�M 2 m@�Cb��ɣL������@� � �M�LɦS�mF���4h� 4d���`F�b0L�`��$ښ�����=A��  �_4���A@V-}�#_�M���a��$U��5F��Z�/�c���������e� kgfyˆvٛ,��rEדd�.�j�܋B @�XI,����]w��w�j�c���_��b�\��K9�W6so'7�����M�)v2��j|��N�O����N��2�껣'�@`����V6������t�/��t������țt�;�pC+����E��	R r��j�Sk������+|͵4���giL:f�yȒӂ�]�{��%r� ����wr\�A.(��q(�4c�4E�4f��,eH�,v\�<���LH�2$|��%�x�N��?���Rj��C@���,, ��I=;�1J
C>hpA�,�N,Qإ6��a�n���Q�4\�i�<"�%-Z�T,�ף��%���Hc��vQ�\b�#yΝV\i�7
&t�#$05��lS�+�qLy�UB)D���2-��^�5()+�]�Q�d��aX`.R��I�c.ռL��gZ@e������Z#���i���;���d��d�ӭ����Q-�E����9e����`ɘ�WPe�d�T*r<���D�r@�1�ū�o9l����#�V�p��
�u��2a� D�P`x��9�;W+���dGXAHϖ2ԩ.��1�ǩ9p���	������1@�i�)z)���o]��h�N����ض3���g�]��BCv�