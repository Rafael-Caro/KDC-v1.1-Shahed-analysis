BZh91AY&SY#Y�� >߀Rx����������`?y���Q�:�.�F-��I �yO4�4�<��j`OB4����a�%	I�jy1S�      A
�z���h��  � �D!)��6�C&4A�DF�� �&L��L �0L�0�D�OD�SlEO���yOOT�=M�b4�.�@���PP�ؠ@M!"IniyR#{�����?s?��i6؂�v�,?i}�X�F� �g��#�������Fm
�{L�o��ۛ�7<�pfb���w�=�����þ�G�,b��Bjrӫ͑����8�l�����k��Z���'�Y2c�~$Q���;i���\��ۛ7!r0�[�$�
i�tC�I�ߒ�rK<p�F���v��1��m�����)�A����D����"a��g�(s�:�j�)�5�#�U��k=zQLٚʱݢw�'JZN��n��hR[�D�5�<����I��Xh cf�s�S�H>�����j�;�5��>z�z��c6�nm�y�d)���S��|�PًD�}�^0���#�Q%Lg��K�HR�҉�v��Ō��2�����-Z�6s�
�WkJℚMJ*;2�92Z�jә����V[r�^<��[���f�q��-�檶�,�X&�6�rSN�����}��)TW:�ș:()�����qX=_v�>~lj��S�՘��!�s������/����6$H�#Y�����7�0�X���=�PG�X�T��
���b�c �@���P����l�&9@_��Q��*Z1H3�i\��ji��U��*!/e��阭�\��jnZ7$��m�������&R�(����Be�ͦ�m@4�hɘjj+�g�B��러���2Gv�Q QԸ��]��o+(l(���	K�#��g�r��ؔ���H�@kۡ�ǣ�����WW������cd��AwU����	��Y�rEF��;�8q��\^N�X�P4eo�n�#o��Q��؍�ⷴ�O�L�f4�Ɔ;ǡ�f츩���V�*-%q�t<��LţCsH%ʋ��ھ�7���G��T�x]"�L(Pb6�*��5u�X�L�L�'b��e��"W�R(E��<AC�2 {arwx�fjȜ��
!)3Ip�J<��Se�@Qd3QC>�bE�O9�CZH�ˁe�Ԗ�W �s�}���`#��0�Z���{M���5���ߡktK�K�^�\�,�W%��/���̶�9�m�'�<�"w'	A��3�$H&��װ��F����௸�d��N�e߷|�NU��S��,��8q���R��Q�\��PUE�%#�>۳Ɯ��q��k�V�.�|�0�t�=qѺ�h_���MnS	R�E����HH�Gh
flM���;�Gb�LJ��,�F%f����n,*X���E�6���Mq�P��.2��<8#��B�vh#o�]��B@�gk�