BZh91AY&SY�ū� =_�Rx����������`<V��.#R��ATCBLI���6�����OSG�OPhf��4�H�S�M�� 2  �h2d�b`ɂd ф``�SS�?Db�4�F��C#C��2d�b`ɂd ф``(	�b&��56��i�e=1@���@�Q(t ��X���B"����N'���������Ѥ�b��j���\�#Q��m3������b��]�F�Dj0`Y��̘�X��$��l�Xa�j�J�jU����;�1���DMq_g�t�'��6���_�ɦ).�A��lhZc@�D*	u
x=�m[��թ<V:!�?bU#M�l�$�X�Zi$�����;w��m�%�5侾��#�㧟��wP�̓|����>���s{���f^��)��e�a����)(�q�40m	�g=U��-�W�����{+��皁q]�T�M��Jq������"l��+8Fp����9�x��m��ړ"�ó���U��}�Tl��>��d�z2��iE�����;E1��dFO-|E�ʴ�5}���B��Ҡ�B���J� ��М��jf�������%�OԿ��p{l\b�u��׌8��ĳ1�By�=�$�A�{�}>�+��1�$z���R,P6�V�k��`Z��
*g��ww�s��x�������}^�gx8�^����	;E��u��|���( ���Wt�ܳ�����9��6�� �)�<��h��;�6ٺ�����9��E����*���c(������C�Z$ĠNrR�)q=��݂/�};�.Nθ�5��t���90eQP��Up}�6��v�M�6�4�a�5V�񳮃 ��\rG^�'NjqHn�8n֙����]�R\a;�M40Fn_�6��� ²F�����&|&j���a0j4�6D D7.�t�r�7��J�d�Q`��B���d���sN))��n0���τd)!zT\�*E�c�m��c����������M���7�̼�8�v���3kGSH#�˿#J� ѳ�\\ �D�^��&$�ab���똲h4X[�4��Rd������4�^\��$XE���;1���.G�� ɚ+���@X�Pʫ%�����ɗ� �,�2������	�yq&��y���fĖ�S�_#��l���"w5���hѤ�j�[�<��%��m/�.�Ť�+��W�S��P;_�ѯ���R���K�3�I�8���3�"T���|K��T�~,ASfJ�]���e�u_��N�>�%���y��|���Ed_r��@!9��(�� �|Ze��I$�mMq�ۋ�^��$a.�:7�o�FE�T�ꁼ̺j�U��B��W`_y����:g��������!Z�m���:��&҅�5�#QRkn�ꛊմT��{��g��r ܏<�����#o�.�p�!��W