BZh91AY&SY))�_ >_�Rx����������`?z۷:E���h �Hm5=�50�i���4h�J=e<�  @�   9�#� �&���0F&�����F!�ѓ@4 4�`�1 �&	�!��L���h�i����z��=TziBz�6�h J�?F(HAa�Z4��i)6�o���8�c�6 �W@�K�GBJ���D���ն"�~r���0�E��Lw�R�ǐ^L�crmXʂ�ڴ*؋^Y�t��Ƌ�g`��c��ɕ��[�-�ͣ�)� 1��5 ��;�2Ґu!�|<�V���K�ͤƔtzY-4*��I �z�+�I&��H^��K������x]���0c�ί���#�`��^Y$Lrϔ�i��aOiy�X��5�iJ�R���R�y_��d$�ݽ:f3���w�We_�2�<���u)"���P�wA�d��+�Tcf,��������S =���_�̶�!kȄ �lQ�"��;\�:�|�6�f�R+�d��fN;JV���M�*(!%XRV�t+eZOl���� ūY�ۦ*�U���F
'Pj�9�L08��2Ȗvh(O��U�f[x8j�S��2;U��Q�a-l�%F��2�x`���%m`��E�?�q�
*�����tP� ~�~'������p/���~��a{�n��*��j�����@}�Aa/��!�!"G�\G�(���o�k糖ܟwSG��_�����Fp��诼y��6Ș�D{9�ٲEƗ�W�~#D�)���$ek��^>��=SbPR�S�9�=�_�0�-ݽG���um���;&�M�0�Q�6��K�ee6+�!�����YZ[x\4�R���.�Z=܉��I!��1+ώ��{ʖ3&]�{ �[B=�ak!���D��*�����ߎ�3�P�u~�����+���� �A�y��N*�vo��%>��9"�#��;��9�ŃQ�þ�� P��)	���I:�1E������!�1��7>����ģ'��,�`K�v=hfUL���Ѥ���6/P��ã�EdP0��FE/ab���砵�UZI�4��Hc���f92�C�%�q��D�P ��9��d��A�p\�*"W��!)����^����0jȳ!��9s�Ӂ�>SC�_B�&��߽%���Ï_������G�P1�z�#^�[+	�'M����m/*]��Iu�]����q�2����vU�w>�}��ԑ<S�������		�������N�z�k U�!eݻ�e���/���OG[]mYMB���V�Չ��EB�0����PJ*�)� {YZ�7(���jMmŷ�/�K˶F�M.լ���H�H9��`bih�R�W�a�#������ɉ���^bGhHܤ[�bb8���$p*^�C5Th\Qp���u͠���uaxϝ�I� �A�h�S���F��]��B@��E|