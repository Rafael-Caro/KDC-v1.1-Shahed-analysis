BZh91AY&SY���? _�Px����߰����P8�h�lư�D�!���)�C��{Tښz#A��j���4��24�#@� M40L�D�I�a4��  ���`LM&L�LM2100	(��ښ��4��� ����H�pd��h"-�ɴ6�l>��BEZK��4��Z��|�{[!�#�)k��C�˪@�/U�-�fx) ��h�l�,[9��+�� P��K	t�>Zp�N�T$�g���Y�e�7��'����N�s}
\�nO��5]	ˇl)�/��9�Q%&�[�!���~W.�394�Y��um�@�}ä�_gI
n�眉�O��b��X�R��M�f�H� ���hh�&*�w,g�#(�h��P��[?U}��U]eW{S��*�2�T��q�
��z��r�B���Ì�Q��KL�̫������opy"!�=�8�S������Xǃ�,���cȑ6�sf�� �i97�)Je���0���-�R�ğ��<5M�������bi��W�
���wyIXiM�r|Z��%�� �y�˴Tgf�^b�|�0:�r�J�9:KT]R�kI��j�:̭�-�tU��j�^�SxS|����Ź�X�0,e��L��iZ�@g�0A��^#"i��!q@<&�0��I)�[�sdo�.�QyEt�,NC�e��m�/W�@]�6p���eB���L۱�dL�|�T�v
*��.�F"�1�V��`�
��A;�~��ĉ"L)6,#�5�܈�̟jb�K��I���5�E��T���Ng%��� `&�p�V�F=YJ^�`Mr��d �2S�.�{�36�d]�rE8P����?