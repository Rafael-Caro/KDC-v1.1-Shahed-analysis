BZh91AY&SY��f� 0_�Rx����������`?zۛ��N�nΝ4h�Hd� &�ڞ��=OP�@2 �&h� i4hL��2��� �`�2��i�"h���0	�	�22 #F9�#� �&���0F&$L��h&54��=G�dz�&S����F�0�@���H,{X�@M!�"Iki|)	&�&�7uzαy� �*��D�~��I\L��HL�b+��@w1{�\�f���D�a�d��g87�T�-�_��;�	��+�E��˶˯����yZ'e����\m뀽����*�!�f���;PמZ��g(<l�P�b��|���i�`���\�A	,������SM�R�I%�������kɊ g(��C��#����z�D Y�oo�{JcZZDK�0��^_B���R�%B �D/ޒx�h���*V�&$�f�¸��C[�T�F��*�5�3'k�ZI��(�e��s�N���?Mc[��@�������K�q,��6� ��C[=��q8�9Œ+Uȑ�j�;[�or�U%�/��U��M�`�L�4�i�IJ�i8
̥V9倢)�F
�o\y2~�91{9b�b�t;���',��_5̠ud8ꏿ�RZ����sq�,��D�����i�7:��m`{]�}zI 5��9*�i����;����Gw3ý�>^[��ګ7������A��}�� >pȻXK��C`BD��n3��c�#m�Ge	䫔)���ߘr����f��]<G�^Q�"c����f�5�L��&f`��1H�����8[�U�R���ְ�`�@�$AB�cK��\�Q�V��n�2\�[�Z\JQ/yU\�NJ�� M�6�t�e�Jq>� �h��W��I�������ؙ�iBƒet/�	%���R�G1�X�zP��4멜�����\����FPS9�����.wd�����"���>NH�H�1N���G�|�
�����
H���a�Se#pe�tF�������0c���>��~82|x�1��1,���C1�f���K����R��ѷ�^B)"P�<�	�P��39<0L��+G�ɓ9!�$Fr�b˄�"K�MD�&"���N�@��p�C ��A:�Yer%|A2��Jij��8�ٙ��}�<W�laP�R�`Ƿ`i#��ʹ�I���a���붃H�#��ٵd#F|��f�Bk#�A������K�b�\H+���������~�>�Fj9Φ�A>a��$O�!(;�jL�	\tf|:����x22W�PJ�sI�'��\����偲dgex��m�X?����DU����NB�S�̆x6��Uؙ�gbb�k�39p�@�DR��y�sIc�I.���|̜KQ��L0Jv+Q皀����}��>i�Q#�Hؤ[qbb2J摸�zf�Dk*\�n�ʦEj�*^�Vk�{o�'���BH�8=�P����1���"�(HP�3c 