BZh91AY&SY$"n _�Px����߰����P8�7Lvͪ�Q"l�=bi��=M��@4 P5I�4�b��  �&�F� $D@I�4������4 �2�101��&$�SF����&�3S#M ����$B
��2����a~�F��M���(H���ګJ�X�����Ii�q��|L���vh����3�B������F�DD��I*MY�o�FR�2�T�o,Y�c�,U���L"_�C��}%(�8���ܾƴ�	�̭X�Y��jɣ2f�p7�;1�7���C�zVf6�����m-_�ݴ�7m�礔n���o��+��a�(n�Lk 9RL��G)K-lF�hk���>i�dN� ��a���*HT5P��>�P�5q(���ZCa	 6����Y��Ǌ'��ȏ2�S>K]	gx\��A�Y���"ڒ�x��O�M��S(��!�Y��[�-�e�B}�M�2����Tb5V�]��ܙ���Hs�����9aF� s�t�,q3��R��������R ��5��O���YB���.�`��$�#O����2��0͘��Tìt�B	W��yV���汩9AT��ꏛdE� ��x�I�0�PM��ʶ���MK�ռ�2Z��e!�F�\��2�ۉ�R�v]6�@�z��b"AQC˓��X�3h>&�� :�kXdU,\W�Ѕ���b7�^b�~Zq�rTP�[2(�\9»x*/1���`ԉ D��`x���h`�҄�S�&���=�}/<ƹ��Y��G�N\Q5� �J����1P�4�V�WW��[FUKo��ع��o�]��B@��M�