BZh91AY&SY�-�� _�Px����߰����P9�ô�Z֌%�6��A��<�h��Ja&b@���� � DD&I�S��(4 ���101��&$�4Ȇ"��OS$���h �OP�*
�ů�Da��46�l:�"��K����ՍnԾ!��C�G�g\q|�k�q�/���3_�z�J��9�����A�`@b"&
-�_[��R�(4<����d���K���<����{q[@����h%��'E�zK�&���K�ՠt2��1��Jg����fci��l��9��������������W�iY!�g��I�	0� �Kٌ����hl;F�h����5�$���0�7��Z�A�`��{��A Ȋ4���zK�Y8oC}p��'��#=D]4|�<��g�\��A�Q���*�Is�i&R�MO��H��!�Y�f c��7�iR�#��^�F�KǮ��/Q˝��竭ݢ4�
5Q��i�L"�;v԰-�K���NJ�;5�Ο97� ��ʻ%�:���E�/�b�\I��W���J��"�蔒��I�t�	汩9��Ut���o"��<��T��
����_�&7o1[�/�� s<�A��=�&!k�y(�(�=��TN˦���T��"�ss$�x\hDX�5��$j�;�HA�j�_�ˊ�� �8�e	�J�����B�+���f^ ��g��oƅ
@��U �n�0ͭ��lF�[:�"��ҥ(y�x+�0|ii�6r�"ui $�h��r�rg�{����벵m�X�~o0���f�2eE��w$S�	��9`