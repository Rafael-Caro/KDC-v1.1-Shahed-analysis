BZh91AY&SY$��@ _�Px����߰����P8�7L�mj��E3$OFj����h i���2yCzH�2m@42�����$DA2����=O#H�� 4���`LM&L�LM2100	)��=��	�S�i���   5�$B
��3����!~�F��M���(H�����J�X�+�K!�����OS-���M�Rwd�7�$���^Q�����c��0�:�I*cwb���6s�*qßo�F��,�|0t�DIC8�JQ��e�-T���֛�R�\�*%��X�qRI�`�~Ҷ�c՚Myt��m;m�3O)�-_���!C���IF��y�xC+�gcFfI�	0� z��
U�=K�����G:qx�U��닧����}1@�$�p��N��%��M�$>�,Ad���?nF�A�ߣL�g(M��2gM�c�cu�������ZVAO�Cؤ�"�CP�� �Q�Д'�u�QT��S�F#Mk���v��<�Ē��;�c��i�:��N�E�&u�`[[�#>��	��&;�هη�PF�J�i>��Fg�ђ@5�Z��u�g�T�lP��-�m�T̒R�1�|�U2�ꥣ�T]1�X�3)~�R{�
�*���V'3p��)�Pȡ�T4�]�}b2N���鵲�U.[
YX�9��#�3D�fr :��͌z9�Խ���l��+g��p��Z.�E/\BǢ�+G8V�Eǝ_�%�bD���G���E\�Bu�sP~�ZH��=�%�I���ʨ��-%����<	���h�ʄjS)["���B�֭�:���k�1�lf�/���ܑN$	?� 