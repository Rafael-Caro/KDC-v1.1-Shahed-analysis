BZh91AY&SY?n� #_�Rx����������`?z۳��7���Δa�a$���1�i�=@4d��4 �$ީ�'�     �A�=$����M�!��� !P��=�F��@4��h��2b10d�2 h�00	#M���?*xS��~�=&!�hi�FL,?d%R
��(HAQ�Z4��@�Z��Z�\�~��%$���F�)�a0F m3�m�����,,h�B��`�\l�٣��0n�k�/��O#C:
�梍�ynw����⴪��1������� �����y@ @<��j`�ҞI:Pg���|8|*�ޭ�&�W	�P_R�e����) R�{�8��Ը���n��j�b-]+�59e`a�~~�m[�L*�7�섉1�����0��(uZv��Y��0�i�v�#C��zЋ�P$#�\�%Xkm�X+�]tLa31������Qg1y�g�yJ�琊��R������e��}1�$��A&�I!��������1��\zH^� ��Y�H�ݾ��,'9fdX�Ί��17x`�D4&H[�c*:T��
LV�Z�����.�&KpB�ZNB:�##��5i��U���@Pͦl�?�R3}�z�����t������YS�AOgW˾��e��əiU�9_<����Bm(X��S��ر\J��)���ڷcO' g�(p� ����`6$H�Sa�x��m�e���=U5�4|r�^9T�?�f��K}#�^��1��x�m��E.��R����SW�H�;�Y6�	��*,xZƪL	�wE[J��(Τ�+�{z'NfM%�TF�v�>�v�`$��(���X��EƛP;6ẸR�O�:�����c�<:I٫	�F���L�iiS2e2^ I.p�	H��._�&P�+A�Ã'}e���	��'k���FP[���� �A��u��o�{�2�i)�[�*8LS��*�߾Z�
-�{���G�נnDb�\�Z�3
�&Z|�[�d�cC���:A��2|x��;�`u������A.5^��e��oyppq�E�xw�1,��J�Fg��ɠ��i&�`l$1Ĉ�@3Y`���IwP�$�1Bt�c�2 ~0������#&5�!��'v�/��P̋�b�F���i�	��X�|�H�۝m���i[��^?��F`z�kP1�j�F[6s[	�N����m.ĺ���AM��^��A�}�Ύ��\�C���pgΒ'�p�Pړ8�D�j�=Y���]�X`uo��b
�A�V%cL�%�
ǰ9-&�k��ЅL&�S��R5{������.3x(��j�����ٍiB������>�[�y,(�j]��4���̊С�b�gI�u��J�=��4����G*����ϥ���&��GpH�R+��1��/�����j�hP�n��JQ�V��U��ݤ����#{�����V"�w$S�	��