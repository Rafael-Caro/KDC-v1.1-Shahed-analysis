BZh91AY&SY��� =߀Rx����������`?z��\��<�@ �L�OT��Sa4j`M1i�=	���BM�l�i @  4� h$��ML�H�m@ 2   �$����MP  4�2dɈ��	�����$H�4M�<��<F��OJx�d��mM����!(;X���@M!�"If��ɀ	\:�����#�e��C��r��`��1�i��"��r���0�����������,n4�=X�������ܳZ���(�\+(j�)ŮW{�I���$����\T�ql�@��C�9�Pb-�{��á���SտP݅.ַ�n��A��#f�8̕@��	�$��w��$��P�&%�}��FC1�͟�����Y�o�|$H{��i3�0��/<�(!��!��L�,h��M;�C��/�W;�Y�ʜ,�:){��$��w���R�(���r�A:]�\4��E�i�Z�]�YP�9���>���lf����m�ϱ&BpP�Ãm�=���d2$N���L�n�-�'u�@ �� R!�I괚FDR�-;�%M����fyVb��Ҡ��K�[# b R�Pb$�IU��?��O"�$K��ȉQ2h���v�#��A/�?"m�r1� ��!�Sm������o�Ō>*��ԋ"�\�����	Lm�ve�R������踐e__�3����	|�B${E���eH��,�h ���������/���[?q�f��z���|�t���G�6�6ȩ��п�f�R���d�S̝;�W��rD:=�{5�Fe�`l7ҹ���uL1-���Kb��̨��V�!.��tM��cM���EYV�8�FwH*���J��D���$7&%9�3_�����^@I-�^b�(C6�ݚ�%v(����큲��x��.3���R1�������$/P�.�W����E	O�}�H�H�1N�ĲG��2	��"�m�@�����	�T��i�����i�c:��C�r�1.d���ˌ	bvǹʉ�Z:��]l��ͫ�GAxtq��� �22.���F���Z�*,�ƚ`j$�%��f92�!�H�𩴒D�\_	�9��d���� �U�W"W��!)���ۯQ�c�M�5dY�����gČP�)��ǯB��۹v������a�_����Y��#�j6pZ׫V�3:BkC��C�6�z]��Iu ��_�O����?9�q��So���lܒ'�p����:�D�j�|v��_��bvs�kY�@ʫ�����d����\����鉾djez��n}������da!u��@E�*))� {MYZ�o�C��jMnŷ�/]�R(�~���]Z�T��2�F���&v��/	�~&<l���LM���<F�"�K��W	J��ب�ʗ.<`4��Z��ʗ�م�?+��A��j=0"�S�ۀ�_�]��BC�#S�