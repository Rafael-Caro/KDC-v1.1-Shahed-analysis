BZh91AY&SYp8�8  �_�Px����߰����P8�0���a(�
b���&&�C#A���% S�����2hh �  ""OIL�O$z��  h�� 挘� ���F	� ���j?S�<=0��@Ѡ� 4h�!AZ5���a~�F��M�W�P�cInj�*�c]�+�C!��������@�Ν�f|�����/��/6�s��L����U��6J�Nc.XMP`����<B�^�7�%�pi|l׼�{a[@�����4���ԝv��Ǽk�R���4�*q,Tq^l(��;�v6������:W���P�DF�IF��xV��aʖP��`�8c&5�-k�a°R���fh?yFZ<
��Q�a��ߤ�u���K��k�F���%�8cs��նY�M\���8�9*����n\���:���ĸ(L~�Kr.�Da�&�\�g�C)6��7�E-^DJŏ�Er
�cU�(O��&T���1�_���s�ٚ$��S���F��F� s�4�X�g����mo�M��R t�l� �L�J�V4���X�(Ac�`e�ŰIc/�F�S�X:)����D�[��Z�� �˅�+R��M��{�H�qB��(%�&$�L��r-. 3��hA��\#"����!r�;�0�=��JTN˦���\�"��`�2m<f��]�D�8d�d�$�5�4����̲���'g-r�]�[�-*Ck��%⨗�	IϧAv'���	���[`��M��ۃ��r'}ڃ��NV+��~t5n�D�$������^8bQq�9	�!E.L�D���,e�/�cb��`_���ܑN$9N 