BZh91AY&SY�2 � >߀Rx����������`?zۜ���r��F�ѐ�B&Й4�S�mL��  h$�10A�h4h ��s F	�0M`�L3JH�if�&��h4�4�& �4d40	�10�"d4�S򧩽L���f���144hɅ�넠�Aq�b�4�D�ť�II����-�u�<�`	�a���_ji+	�0�i�؊���K��Ƌ�5j����K(�.S蟆��3)3n6oµ������	Y�|�B�Q������NgV���TX46�G��F�9�X�j�f�*� ?N���o�H�U�;I�Pi�y-v0�)�i�[��p���.��s�g�/�c9o���o�Fs`���\�&9m"{�0��T���Kb�F��MT�:]��	g0��]�hEq�#��$,)��2��7�Rt�i�L�Yu��H*��3�0�H"L��
YЬZP���J��Tv7��u��]mĈA  \͊:".?/w��L�9ѡ�W����El%ʯ�嬢�&ls���^�V$a���c<�QM�����C�8�/T��wCx!,�4|zD��rb�r��f˝ޚG��Y׎�|��@�˦,�1����pFiI,���Eqv�%u��Xz$l"Ϡ+����l�Kd���aNi���x"B�;��.͌yyn���y��
-�W�����.�	v��6$H��1ٞ<Q�6�;� �J�B�>�v�V��?�N[ 2ÜY����-lg=����1���4L�����@������n�W���|��lJ,���ρ�9}�"������n[U�r�k��F�L���w���t�W�0Cmb:VW�\TJ�i�#ү����G-*�@������&h�P��L���	%���NdG1���a�B�"�H�pW��r��&VΏ��)XAL�k$H2^�r�%]�7�D��|���pH�1N��\�׾��R��ɉ�|#sհ.4-A���n#�.�r?fzƘ���Sc�y��x2|x��M��:Gq�g�f�- ���A�x ѷ��88�Q���yr�L��38�PL�j+W�ɦbI�"Y�a��	D�*��$LE���`���ጆ@�-��U
��b%l!2��Jij��8��{PA�1H��ي��H�-nҭ�H�7�4�&7S<�.?3����?"G6�cfՐ��j11�&�8k6�/nᴾĺ�;Iq �Ғ^��FqA���m�E�s�M^b|�N��<����ԙ��\{3::�{H�M�쌕�F�Ĕ�1�lUU�
�eF��j�h���6��K��qqMx�x5S�Ёu��!��k�Tڜ�9�,�l�39o�$�����^沶D�H�]�ct��
�Mf�1ƥ(<��z�9�k���$lR.�\LFC�[�n(Z�J�1*X�n�ʦEj��-k��F{��OyT9��9ȡa/%[�.�p�!�dA`