BZh91AY&SY���% 0߀Rx����������`?z���ִ�a�gOMe��d�SژҞL$ڞ����@ �&F�H�54i�F�S&���bOQI�CG�42  �4  a ��m@ 4@ @ � �`�2��H�2&�M)�S�6�����D���4����Pu����@��B"R���H��Z=����!�����	��@{B� ��#!��m3�m��_�����������@$@3e��wo�SD�\�����mZ|"מ/,��T����R��G)����&�0$����W!B!�&s��vsa��F#Q�������wq��kt�mZ�rh�p���H���#q$��99{#����PFkj�l��,0��k�?�V�*l��䔊F6��=C��u���&�h���C��d�s���� �:bfI^N��&b3t��kba`h�J��#�Qñp�0�<`�`5��M�~��ޯ�	^��˫�x�����7��=	2��w�K1p�\֖��� ����7���	C��h`�_�"�x�e���d�4E4��\,��,�V*�a�Q�1|��O �Ũ�W:���tN=��N_z�U��]	�eݑ�]r�����2G[.�/�Fl&��v�[X"������ ��+��P7�$�dO���
���.Z�Tße�r��c��aU��+z{A��>pȻP`%�����;���y��z?�f��Q�=�ۡQ+L��p3��Fm��篴zE��L�TG~��:$���
�/�h��E��^.3�kl�b�Q�m`Nl���L�s"�.Y+5��I�f�7g26�����n�����b{7Y])64ڀi�4U��4�pg)��~���#è���q ��dW~�i�604�-�w�)t�l�JDG1�X���4W$f8)�3+��c�q��~߂�+��+��1�B	��.wnV߃{`4IRi�NNQ�I���#˾���b�É��ࡒ:��E�?eM��c��*�y��`B�cC�o��u��.e8�M7���<Z���Z8�A<p^�� ѳ�^B+%�0�
<�$Ha~XA%��dɁ���$��2�˄�"W;�PE�𝠁��ጆ@�-n�v3r&�:%#&h�Eר�1�ј��@��0b����)c�U�hi#����I��������K 6�62p�1�Z�cZ�33��-��g�Kȗ ��\H-���}�q�Pz�a�_#�R�GaNa��$S$�!(;�bL�	�\ud|;L<���LU�F���	A��A��xD�R4P}B�"�-`-w�j�.,)"o�D�t YE=<�g�h+i_=��s:�S-4fg-��x�E./3��}q%yy`�f�鑄���b`%�	�y� T�h��d4ט��I�I���7ű�iR��*��X�m�����m
��׍�>7ꗼ��B�pm"�u��_���)�%�i(