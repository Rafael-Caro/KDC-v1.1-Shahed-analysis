BZh91AY&SY��A" 0߀Rx����������`?zۜ�Y��t
5 F��Jz�F�j~�h����4� 4D���H��4�����0L@0	�h�h`ba��IC�4�ѩ���yA��F�h@� �`�2��H�&�&��'��ڞDf�5=OQ�hd4dʂ�As��i.!KcK��$��?��ky" BRF�(%���%B`��"@�g��l�y�����E��- � ��*�e�0�z8��[ �2.E���������Kw�+T���7�֒� X71���6R���i����uhSW\6����ro�QԴ�_̂�(��}�I$
z�]�d�K}m��sK�=z�0�^��d#H�~I���~�2��鄉��m"A�{�v�2�y)!M��D/�7"���npQMA�
�Ƥ�(2Y)ITd��j��-5j��MָgKҷ���⚻�k���N+�ӑ.�a@���0 � N(���2��F�U�`��A#@���Ui���tU�u����RQ|a� �n�R��c$��45�<"*���n��I�&W���
>[se�����|[>��Iu�_j�f�s��B��T�۔ݪ�]��fy��"d`��gd�lgwQ����oGפ eS�-�Ч<�~<��#�����c�۲_UƩ��m�XUn �oOh3���]�.%������o4�cڏ����Qzy�g
h�-r�b9\ӯ��o��_��rȘ��;��l�cf��!�f,�,R�N4��'|��}#�z&Ġ�&��9�=�Lp��ޭ�u�ܹj��,��/��n��8�0���8���+9�cM���F��N'��2��~��G?	�e ���..����,\_���w!9��K��$�I\��p�ꅯ�l'W��R2�5tc$H3^quS5n{��T����}.H�H�1N�ȺG_<���G&�
�ۡ1�a�Sh#ta��'Zd}�+��0c���>�`}�d��&�����b����8A.7]��E��wY�pq��!�H�S.1ο=�����&4�A!�$F��ie�"K��!$���A�'h `�8c!��k����f]Q���	Hd�4�)���%6b� ��H%��Mୂ
V�l�,$wGhƪ�[/]3���g���`x�;�����b5h��l6VY�9M�[��_R]!����[qY/u�H��?1�oI�\�c��O�5��%hnI��H�\��E��y�a�T����d
Y���sI�'委�NJ��Fّ������29�b��SE .��T�񉒒�����c��������ZU��q�Ľ"Im��ֻ�̝��H�[�%�"�T�7�FrXT��^���XM�5�H�	T��.LFc�ldo*`�a�U[��gc2�m�pk�{��'�A��R9\=d����A��ܑN$$�PH�