BZh91AY&SY��� #_�Rx����������`?z������u�C��QS�2���I��z� 䆞�1 ! M$�L� 22 � ����@�A���!���  �(�S�'��O@G�m!�4���8ɓ&# &L �# C �"d����I��=O� �h6�LLn?�����	� ��I-�/
��������_��6 �W�t��N�b1�?�؊����/��h�F@,@8Յ�ƞ�u�һik�*��P}��ɪd�h�K��h�Ǔlo���� ^L�?3�Ea 2�e�"�'<�ʰ�J�̈́*���������h>�7Sn/�.��$Ih�G�I�<�Y�i���i�d��((`��r���X���
C����H%�a �:���r�4J"C��9� ţ�:m��T���ȹ���%iv���1�̶ia;_+ө��.qP��
F��eꙢ�"4n�g�>gy�b9�  ��tDY�sz�j�7���p/iK8�h"��⫂�=U�U�V�K�+iу#E`�&Q �f0RN�cD;�1Q��TiPa�_%թ�s� lӌ-*�*�\f��.�7,$֛CS53?ys4���4	�Rd:�(���Iӭ��a��wW�#�� 4�����x�cC�:8�#���tWe�Q��J6��X��n�g���]�,%��0$w3A���}M�]�w���p����_+r���槬y�R&>X��sm��T�|3/���$��	�!�₧�$�G���}��Ө	P���';�y�)*�MN�glQ�����#�t��}�R��H耪Y�r�d�V�0CӦ��*ԧ�ΙCV8�i]:���$p�BW�bSv|i���,dL�������-b�3Z�3A$���6��2�g���:?g�H��j
h<�l�A �yE���wY�HR(J}��rE�F��v%�:�Aۙ��ڷMt����8j��>ދk��G��è�'�yr�1�����}ܠ�x�2}���X�ñ�C4�3��y����j5�8z��{�E$\Xc#Iu�,Xb2:��SAeE�Li��I�"Zc��	D�
��$LE��`���ጆ@�.7A
�Yer%|�2��Jik��q)��,�2x�E;��ZUD@�!��"�W�+��/s%�	�����q#��lڳ�F�f�e!5���ۼ����K�4��Av�����E��8�L(�:������D�N��6�ΈH�MRnG��_�.19�j5- ��UrW4ӚL�=_�y(��:�8-�G���o���<��3"���@W�\��a�F2��M
���X��TDS�7}�$����=s�����L�p�D�p16Z8�^J�L0$v�?WL�X��k�H�8ԋr&#1Ԯ9
��d���K�'$u3+V�YR����g���{�:bkG�� At{�[�.�p�!!O�.